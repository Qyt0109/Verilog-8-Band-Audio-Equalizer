module filter (
    // system signal ports
    input clk,
    input clk_enable,
    input rst,

    // filter module ports
    input signed [15:0] filter_in,  // signed integer 16. [-32768, 32768 - 1]

    output signed [15:0] filter_out  // signed integer 16. [-32768, 32768 - 1]
);
  // region coeffs
  // Store the coefficients internally
  localparam NUMBER_OF_TAPS = 63;
  parameter signed [15:0] coeffs[0:NUMBER_OF_TAPS-1] = {
    16'b1111111111110110,
    16'b1111111111100001,
    16'b1111111111001011,
    16'b1111111110111000,
    16'b1111111110101001,
    16'b1111111110100111,
    16'b1111111110110111,
    16'b1111111111100001,
    16'b0000000000100110,
    16'b0000000010000011,
    16'b0000000011101011,
    16'b0000000101001010,
    16'b0000000110000111,
    16'b0000000110000111,
    16'b0000000100110010,
    16'b0000000001111101,
    16'b1111111101101111,
    16'b1111111000100001,
    16'b1111110011000101,
    16'b1111101110011001,
    16'b1111101011101011,
    16'b1111101100000101,
    16'b1111110000100011,
    16'b1111111001101011,
    16'b0000000111011101,
    16'b0000011001010101,
    16'b0000101110000101,
    16'b0001000011111111,
    16'b0001011001000010,
    16'b0001101011001001,
    16'b0001111000011011,
    16'b0001111111011100,
    16'b0001111111011100,
    16'b0001111000011011,
    16'b0001101011001001,
    16'b0001011001000010,
    16'b0001000011111111,
    16'b0000101110000101,
    16'b0000011001010101,
    16'b0000000111011101,
    16'b1111111001101011,
    16'b1111110000100011,
    16'b1111101100000101,
    16'b1111101011101011,
    16'b1111101110011001,
    16'b1111110011000101,
    16'b1111111000100001,
    16'b1111111101101111,
    16'b0000000001111101,
    16'b0000000100110010,
    16'b0000000110000111,
    16'b0000000110000111,
    16'b0000000101001010,
    16'b0000000011101011,
    16'b0000000010000011,
    16'b0000000000100110,
    16'b1111111111100001,
    16'b1111111110110111,
    16'b1111111110100111,
    16'b1111111110101001,
    16'b1111111110111000,
    16'b1111111111001011,
    16'b1111111111100001,
    16'b1111111111110110
  };
  // endregion coeffs

  // region counter
  wire [5:0] current_count;

  counter counter_inst (
      .clk(clk),
      .clk_enable(clk_enable),
      .rst(rst),

      .current_count(current_count)
  );
  // endregion counter



endmodule
