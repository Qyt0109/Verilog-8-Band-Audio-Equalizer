// python compile.py filter counter.v phase_check.v delay_pipeline.v input_register.v write_done_capture.v coeffs_control.v compute.v filter_impluse_tb.v filter.v
`timescale 1 ns / 1 ns

module filter_impluse_tb;

  // Function definitions
  function signed [15:0] abs;
    input signed [15:0] arg;
    begin
      abs = arg > 0 ? arg : -arg;
    end
  endfunction  // function abs

  task filter_in_data_log_task;
    input clk;
    input reset;
    input rdenb;
    inout [7:0] addr;
    output done;
    begin

      // Counter to generate the address
      if (reset == 1) addr = 0;
      else begin
        if (rdenb == 1) begin
          if (addr == 129) addr = addr;
          else addr = addr + 1;
        end
      end

      // Done Signal generation.
      if (reset == 1) done = 0;
      else if (addr == 129) done = 1;
      else done = 0;

    end
  endtask  // filter_in_data_log_task

  task write_enable_data_log_task;
    input clk;
    input reset;
    input rdenb;
    inout [13:0] addr;
    output done;
    begin

      // Counter to generate the address
      if (reset == 1) addr = 0;
      else begin
        if (rdenb == 1) begin
          if (addr == 8319) addr = addr;
          else addr = addr + 1;
        end
      end

      // Done Signal generation.
      if (reset == 1) done = 0;
      else if (addr == 8319) done = 1;
      else done = 0;

    end
  endtask  // write_enable_data_log_task

  task write_done_data_log_task;
    input clk;
    input reset;
    input rdenb;
    inout [13:0] addr;
    output done;
    begin

      // Counter to generate the address
      if (reset == 1) addr = 0;
      else begin
        if (rdenb == 1) begin
          if (addr == 8319) addr = addr;
          else addr = addr + 1;
        end
      end

      // Done Signal generation.
      if (reset == 1) done = 0;
      else if (addr == 8319) done = 1;
      else done = 0;

    end
  endtask  // write_done_data_log_task

  task write_address_data_log_task;
    input clk;
    input reset;
    input rdenb;
    inout [13:0] addr;
    output done;
    begin

      // Counter to generate the address
      if (reset == 1) addr = 0;
      else begin
        if (rdenb == 1) begin
          if (addr == 8319) addr = addr;
          else addr = addr + 1;
        end
      end

      // Done Signal generation.
      if (reset == 1) done = 0;
      else if (addr == 8319) done = 1;
      else done = 0;

    end
  endtask  // write_address_data_log_task

  task coeffs_in_data_log_task;
    input clk;
    input reset;
    input rdenb;
    inout [13:0] addr;
    output done;
    begin

      // Counter to generate the address
      if (reset == 1) addr = 0;
      else begin
        if (rdenb == 1) begin
          if (addr == 8319) addr = addr;
          else addr = addr + 1;
        end
      end

      // Done Signal generation.
      if (reset == 1) done = 0;
      else if (addr == 8319) done = 1;
      else done = 0;

    end
  endtask  // coeffs_in_data_log_task

  task filter_out_task;
    input clk;
    input reset;
    input rdenb;
    inout [7:0] addr;
    output done;
    begin

      // Counter to generate the address
      if (reset == 1) addr = 0;
      else begin
        if (rdenb == 1) begin
          if (addr == 129) addr = addr;
          else addr = #1 addr + 1;
        end
      end

      // Done Signal generation.
      if (reset == 1) done = 0;
      else if (addr == 129) done = 1;
      else done = 0;

    end
  endtask  // filter_out_task

  // Constants
  parameter clk_high = 5;
  parameter clk_low = 5;
  parameter clk_period = 10;
  parameter clk_hold = 2;

  reg signed [15:0] filter_in_data_log_force[0:129];
  reg write_enable_data_log_force[0:8319];
  reg write_done_data_log_force[0:8319];
  reg [5:0] write_address_data_log_force[0:8319];
  reg signed [15:0] coeffs_in_data_log_force[0:8319];
  reg signed [15:0] filter_out_expected[0:129];


  // **************************************
  initial  //Input & Output data
    begin
      $dumpfile("./Simulate/impulse.vcd");
      $dumpvars;
      // Input data for filter_in_data_log
      filter_in_data_log_force[  0] <= 16'h0000;
      filter_in_data_log_force[  1] <= 16'h0000;
      filter_in_data_log_force[  2] <= 16'h7fff;
      filter_in_data_log_force[  3] <= 16'h0000;
      filter_in_data_log_force[  4] <= 16'h0000;
      filter_in_data_log_force[  5] <= 16'h0000;
      filter_in_data_log_force[  6] <= 16'h0000;
      filter_in_data_log_force[  7] <= 16'h0000;
      filter_in_data_log_force[  8] <= 16'h0000;
      filter_in_data_log_force[  9] <= 16'h0000;
      filter_in_data_log_force[ 10] <= 16'h0000;
      filter_in_data_log_force[ 11] <= 16'h0000;
      filter_in_data_log_force[ 12] <= 16'h0000;
      filter_in_data_log_force[ 13] <= 16'h0000;
      filter_in_data_log_force[ 14] <= 16'h0000;
      filter_in_data_log_force[ 15] <= 16'h0000;
      filter_in_data_log_force[ 16] <= 16'h0000;
      filter_in_data_log_force[ 17] <= 16'h0000;
      filter_in_data_log_force[ 18] <= 16'h0000;
      filter_in_data_log_force[ 19] <= 16'h0000;
      filter_in_data_log_force[ 20] <= 16'h0000;
      filter_in_data_log_force[ 21] <= 16'h0000;
      filter_in_data_log_force[ 22] <= 16'h0000;
      filter_in_data_log_force[ 23] <= 16'h0000;
      filter_in_data_log_force[ 24] <= 16'h0000;
      filter_in_data_log_force[ 25] <= 16'h0000;
      filter_in_data_log_force[ 26] <= 16'h0000;
      filter_in_data_log_force[ 27] <= 16'h0000;
      filter_in_data_log_force[ 28] <= 16'h0000;
      filter_in_data_log_force[ 29] <= 16'h0000;
      filter_in_data_log_force[ 30] <= 16'h0000;
      filter_in_data_log_force[ 31] <= 16'h0000;
      filter_in_data_log_force[ 32] <= 16'h0000;
      filter_in_data_log_force[ 33] <= 16'h0000;
      filter_in_data_log_force[ 34] <= 16'h0000;
      filter_in_data_log_force[ 35] <= 16'h0000;
      filter_in_data_log_force[ 36] <= 16'h0000;
      filter_in_data_log_force[ 37] <= 16'h0000;
      filter_in_data_log_force[ 38] <= 16'h0000;
      filter_in_data_log_force[ 39] <= 16'h0000;
      filter_in_data_log_force[ 40] <= 16'h0000;
      filter_in_data_log_force[ 41] <= 16'h0000;
      filter_in_data_log_force[ 42] <= 16'h0000;
      filter_in_data_log_force[ 43] <= 16'h0000;
      filter_in_data_log_force[ 44] <= 16'h0000;
      filter_in_data_log_force[ 45] <= 16'h0000;
      filter_in_data_log_force[ 46] <= 16'h0000;
      filter_in_data_log_force[ 47] <= 16'h0000;
      filter_in_data_log_force[ 48] <= 16'h0000;
      filter_in_data_log_force[ 49] <= 16'h0000;
      filter_in_data_log_force[ 50] <= 16'h0000;
      filter_in_data_log_force[ 51] <= 16'h0000;
      filter_in_data_log_force[ 52] <= 16'h0000;
      filter_in_data_log_force[ 53] <= 16'h0000;
      filter_in_data_log_force[ 54] <= 16'h0000;
      filter_in_data_log_force[ 55] <= 16'h0000;
      filter_in_data_log_force[ 56] <= 16'h0000;
      filter_in_data_log_force[ 57] <= 16'h0000;
      filter_in_data_log_force[ 58] <= 16'h0000;
      filter_in_data_log_force[ 59] <= 16'h0000;
      filter_in_data_log_force[ 60] <= 16'h0000;
      filter_in_data_log_force[ 61] <= 16'h0000;
      filter_in_data_log_force[ 62] <= 16'h0000;
      filter_in_data_log_force[ 63] <= 16'h0000;
      filter_in_data_log_force[ 64] <= 16'h0000;
      filter_in_data_log_force[ 65] <= 16'h0000;
      filter_in_data_log_force[ 66] <= 16'h0000;
      filter_in_data_log_force[ 67] <= 16'h0000;
      filter_in_data_log_force[ 68] <= 16'h0000;
      filter_in_data_log_force[ 69] <= 16'h0000;
      filter_in_data_log_force[ 70] <= 16'h0000;
      filter_in_data_log_force[ 71] <= 16'h0000;
      filter_in_data_log_force[ 72] <= 16'h0000;
      filter_in_data_log_force[ 73] <= 16'h0000;
      filter_in_data_log_force[ 74] <= 16'h0000;
      filter_in_data_log_force[ 75] <= 16'h0000;
      filter_in_data_log_force[ 76] <= 16'h0000;
      filter_in_data_log_force[ 77] <= 16'h0000;
      filter_in_data_log_force[ 78] <= 16'h0000;
      filter_in_data_log_force[ 79] <= 16'h0000;
      filter_in_data_log_force[ 80] <= 16'h0000;
      filter_in_data_log_force[ 81] <= 16'h0000;
      filter_in_data_log_force[ 82] <= 16'h7fff;
      filter_in_data_log_force[ 83] <= 16'h7fff;
      filter_in_data_log_force[ 84] <= 16'h7fff;
      filter_in_data_log_force[ 85] <= 16'h7fff;
      filter_in_data_log_force[ 86] <= 16'h7fff;
      filter_in_data_log_force[ 87] <= 16'h7fff;
      filter_in_data_log_force[ 88] <= 16'h7fff;
      filter_in_data_log_force[ 89] <= 16'h7fff;
      filter_in_data_log_force[ 90] <= 16'h7fff;
      filter_in_data_log_force[ 91] <= 16'h7fff;
      filter_in_data_log_force[ 92] <= 16'h7fff;
      filter_in_data_log_force[ 93] <= 16'h7fff;
      filter_in_data_log_force[ 94] <= 16'h7fff;
      filter_in_data_log_force[ 95] <= 16'h7fff;
      filter_in_data_log_force[ 96] <= 16'h7fff;
      filter_in_data_log_force[ 97] <= 16'h7fff;
      filter_in_data_log_force[ 98] <= 16'h7fff;
      filter_in_data_log_force[ 99] <= 16'h7fff;
      filter_in_data_log_force[100] <= 16'h7fff;
      filter_in_data_log_force[101] <= 16'h7fff;
      filter_in_data_log_force[102] <= 16'h7fff;
      filter_in_data_log_force[103] <= 16'h7fff;
      filter_in_data_log_force[104] <= 16'h7fff;
      filter_in_data_log_force[105] <= 16'h7fff;
      filter_in_data_log_force[106] <= 16'h7fff;
      filter_in_data_log_force[107] <= 16'h7fff;
      filter_in_data_log_force[108] <= 16'h7fff;
      filter_in_data_log_force[109] <= 16'h7fff;
      filter_in_data_log_force[110] <= 16'h7fff;
      filter_in_data_log_force[111] <= 16'h7fff;
      filter_in_data_log_force[112] <= 16'h7fff;
      filter_in_data_log_force[113] <= 16'h7fff;
      filter_in_data_log_force[114] <= 16'h7fff;
      filter_in_data_log_force[115] <= 16'h7fff;
      filter_in_data_log_force[116] <= 16'h7fff;
      filter_in_data_log_force[117] <= 16'h7fff;
      filter_in_data_log_force[118] <= 16'h7fff;
      filter_in_data_log_force[119] <= 16'h7fff;
      filter_in_data_log_force[120] <= 16'h7fff;
      filter_in_data_log_force[121] <= 16'h7fff;
      filter_in_data_log_force[122] <= 16'h7fff;
      filter_in_data_log_force[123] <= 16'h7fff;
      filter_in_data_log_force[124] <= 16'h7fff;
      filter_in_data_log_force[125] <= 16'h7fff;
      filter_in_data_log_force[126] <= 16'h7fff;
      filter_in_data_log_force[127] <= 16'h7fff;
      filter_in_data_log_force[128] <= 16'h7fff;
      filter_in_data_log_force[129] <= 16'h7fff;

      // Input data for write_enable_data_log
      write_enable_data_log_force[   0] <= 1'h1;
      write_enable_data_log_force[   1] <= 1'h1;
      write_enable_data_log_force[   2] <= 1'h1;
      write_enable_data_log_force[   3] <= 1'h1;
      write_enable_data_log_force[   4] <= 1'h1;
      write_enable_data_log_force[   5] <= 1'h1;
      write_enable_data_log_force[   6] <= 1'h1;
      write_enable_data_log_force[   7] <= 1'h1;
      write_enable_data_log_force[   8] <= 1'h1;
      write_enable_data_log_force[   9] <= 1'h1;
      write_enable_data_log_force[  10] <= 1'h1;
      write_enable_data_log_force[  11] <= 1'h1;
      write_enable_data_log_force[  12] <= 1'h1;
      write_enable_data_log_force[  13] <= 1'h1;
      write_enable_data_log_force[  14] <= 1'h1;
      write_enable_data_log_force[  15] <= 1'h1;
      write_enable_data_log_force[  16] <= 1'h1;
      write_enable_data_log_force[  17] <= 1'h1;
      write_enable_data_log_force[  18] <= 1'h1;
      write_enable_data_log_force[  19] <= 1'h1;
      write_enable_data_log_force[  20] <= 1'h1;
      write_enable_data_log_force[  21] <= 1'h1;
      write_enable_data_log_force[  22] <= 1'h1;
      write_enable_data_log_force[  23] <= 1'h1;
      write_enable_data_log_force[  24] <= 1'h1;
      write_enable_data_log_force[  25] <= 1'h1;
      write_enable_data_log_force[  26] <= 1'h1;
      write_enable_data_log_force[  27] <= 1'h1;
      write_enable_data_log_force[  28] <= 1'h1;
      write_enable_data_log_force[  29] <= 1'h1;
      write_enable_data_log_force[  30] <= 1'h1;
      write_enable_data_log_force[  31] <= 1'h1;
      write_enable_data_log_force[  32] <= 1'h1;
      write_enable_data_log_force[  33] <= 1'h1;
      write_enable_data_log_force[  34] <= 1'h1;
      write_enable_data_log_force[  35] <= 1'h1;
      write_enable_data_log_force[  36] <= 1'h1;
      write_enable_data_log_force[  37] <= 1'h1;
      write_enable_data_log_force[  38] <= 1'h1;
      write_enable_data_log_force[  39] <= 1'h1;
      write_enable_data_log_force[  40] <= 1'h1;
      write_enable_data_log_force[  41] <= 1'h1;
      write_enable_data_log_force[  42] <= 1'h1;
      write_enable_data_log_force[  43] <= 1'h1;
      write_enable_data_log_force[  44] <= 1'h1;
      write_enable_data_log_force[  45] <= 1'h1;
      write_enable_data_log_force[  46] <= 1'h1;
      write_enable_data_log_force[  47] <= 1'h1;
      write_enable_data_log_force[  48] <= 1'h1;
      write_enable_data_log_force[  49] <= 1'h1;
      write_enable_data_log_force[  50] <= 1'h1;
      write_enable_data_log_force[  51] <= 1'h1;
      write_enable_data_log_force[  52] <= 1'h1;
      write_enable_data_log_force[  53] <= 1'h1;
      write_enable_data_log_force[  54] <= 1'h1;
      write_enable_data_log_force[  55] <= 1'h1;
      write_enable_data_log_force[  56] <= 1'h1;
      write_enable_data_log_force[  57] <= 1'h1;
      write_enable_data_log_force[  58] <= 1'h1;
      write_enable_data_log_force[  59] <= 1'h1;
      write_enable_data_log_force[  60] <= 1'h1;
      write_enable_data_log_force[  61] <= 1'h1;
      write_enable_data_log_force[  62] <= 1'h1;
      write_enable_data_log_force[  63] <= 1'h1;
      write_enable_data_log_force[  64] <= 1'h0;
      write_enable_data_log_force[  65] <= 1'h0;
      write_enable_data_log_force[  66] <= 1'h0;
      write_enable_data_log_force[  67] <= 1'h0;
      write_enable_data_log_force[  68] <= 1'h0;
      write_enable_data_log_force[  69] <= 1'h0;
      write_enable_data_log_force[  70] <= 1'h0;
      write_enable_data_log_force[  71] <= 1'h0;
      write_enable_data_log_force[  72] <= 1'h0;
      write_enable_data_log_force[  73] <= 1'h0;
      write_enable_data_log_force[  74] <= 1'h0;
      write_enable_data_log_force[  75] <= 1'h0;
      write_enable_data_log_force[  76] <= 1'h0;
      write_enable_data_log_force[  77] <= 1'h0;
      write_enable_data_log_force[  78] <= 1'h0;
      write_enable_data_log_force[  79] <= 1'h0;
      write_enable_data_log_force[  80] <= 1'h0;
      write_enable_data_log_force[  81] <= 1'h0;
      write_enable_data_log_force[  82] <= 1'h0;
      write_enable_data_log_force[  83] <= 1'h0;
      write_enable_data_log_force[  84] <= 1'h0;
      write_enable_data_log_force[  85] <= 1'h0;
      write_enable_data_log_force[  86] <= 1'h0;
      write_enable_data_log_force[  87] <= 1'h0;
      write_enable_data_log_force[  88] <= 1'h0;
      write_enable_data_log_force[  89] <= 1'h0;
      write_enable_data_log_force[  90] <= 1'h0;
      write_enable_data_log_force[  91] <= 1'h0;
      write_enable_data_log_force[  92] <= 1'h0;
      write_enable_data_log_force[  93] <= 1'h0;
      write_enable_data_log_force[  94] <= 1'h0;
      write_enable_data_log_force[  95] <= 1'h0;
      write_enable_data_log_force[  96] <= 1'h0;
      write_enable_data_log_force[  97] <= 1'h0;
      write_enable_data_log_force[  98] <= 1'h0;
      write_enable_data_log_force[  99] <= 1'h0;
      write_enable_data_log_force[ 100] <= 1'h0;
      write_enable_data_log_force[ 101] <= 1'h0;
      write_enable_data_log_force[ 102] <= 1'h0;
      write_enable_data_log_force[ 103] <= 1'h0;
      write_enable_data_log_force[ 104] <= 1'h0;
      write_enable_data_log_force[ 105] <= 1'h0;
      write_enable_data_log_force[ 106] <= 1'h0;
      write_enable_data_log_force[ 107] <= 1'h0;
      write_enable_data_log_force[ 108] <= 1'h0;
      write_enable_data_log_force[ 109] <= 1'h0;
      write_enable_data_log_force[ 110] <= 1'h0;
      write_enable_data_log_force[ 111] <= 1'h0;
      write_enable_data_log_force[ 112] <= 1'h0;
      write_enable_data_log_force[ 113] <= 1'h0;
      write_enable_data_log_force[ 114] <= 1'h0;
      write_enable_data_log_force[ 115] <= 1'h0;
      write_enable_data_log_force[ 116] <= 1'h0;
      write_enable_data_log_force[ 117] <= 1'h0;
      write_enable_data_log_force[ 118] <= 1'h0;
      write_enable_data_log_force[ 119] <= 1'h0;
      write_enable_data_log_force[ 120] <= 1'h0;
      write_enable_data_log_force[ 121] <= 1'h0;
      write_enable_data_log_force[ 122] <= 1'h0;
      write_enable_data_log_force[ 123] <= 1'h0;
      write_enable_data_log_force[ 124] <= 1'h0;
      write_enable_data_log_force[ 125] <= 1'h0;
      write_enable_data_log_force[ 126] <= 1'h0;
      write_enable_data_log_force[ 127] <= 1'h0;
      write_enable_data_log_force[ 128] <= 1'h0;
      write_enable_data_log_force[ 129] <= 1'h0;
      write_enable_data_log_force[ 130] <= 1'h0;
      write_enable_data_log_force[ 131] <= 1'h0;
      write_enable_data_log_force[ 132] <= 1'h0;
      write_enable_data_log_force[ 133] <= 1'h0;
      write_enable_data_log_force[ 134] <= 1'h0;
      write_enable_data_log_force[ 135] <= 1'h0;
      write_enable_data_log_force[ 136] <= 1'h0;
      write_enable_data_log_force[ 137] <= 1'h0;
      write_enable_data_log_force[ 138] <= 1'h0;
      write_enable_data_log_force[ 139] <= 1'h0;
      write_enable_data_log_force[ 140] <= 1'h0;
      write_enable_data_log_force[ 141] <= 1'h0;
      write_enable_data_log_force[ 142] <= 1'h0;
      write_enable_data_log_force[ 143] <= 1'h0;
      write_enable_data_log_force[ 144] <= 1'h0;
      write_enable_data_log_force[ 145] <= 1'h0;
      write_enable_data_log_force[ 146] <= 1'h0;
      write_enable_data_log_force[ 147] <= 1'h0;
      write_enable_data_log_force[ 148] <= 1'h0;
      write_enable_data_log_force[ 149] <= 1'h0;
      write_enable_data_log_force[ 150] <= 1'h0;
      write_enable_data_log_force[ 151] <= 1'h0;
      write_enable_data_log_force[ 152] <= 1'h0;
      write_enable_data_log_force[ 153] <= 1'h0;
      write_enable_data_log_force[ 154] <= 1'h0;
      write_enable_data_log_force[ 155] <= 1'h0;
      write_enable_data_log_force[ 156] <= 1'h0;
      write_enable_data_log_force[ 157] <= 1'h0;
      write_enable_data_log_force[ 158] <= 1'h0;
      write_enable_data_log_force[ 159] <= 1'h0;
      write_enable_data_log_force[ 160] <= 1'h0;
      write_enable_data_log_force[ 161] <= 1'h0;
      write_enable_data_log_force[ 162] <= 1'h0;
      write_enable_data_log_force[ 163] <= 1'h0;
      write_enable_data_log_force[ 164] <= 1'h0;
      write_enable_data_log_force[ 165] <= 1'h0;
      write_enable_data_log_force[ 166] <= 1'h0;
      write_enable_data_log_force[ 167] <= 1'h0;
      write_enable_data_log_force[ 168] <= 1'h0;
      write_enable_data_log_force[ 169] <= 1'h0;
      write_enable_data_log_force[ 170] <= 1'h0;
      write_enable_data_log_force[ 171] <= 1'h0;
      write_enable_data_log_force[ 172] <= 1'h0;
      write_enable_data_log_force[ 173] <= 1'h0;
      write_enable_data_log_force[ 174] <= 1'h0;
      write_enable_data_log_force[ 175] <= 1'h0;
      write_enable_data_log_force[ 176] <= 1'h0;
      write_enable_data_log_force[ 177] <= 1'h0;
      write_enable_data_log_force[ 178] <= 1'h0;
      write_enable_data_log_force[ 179] <= 1'h0;
      write_enable_data_log_force[ 180] <= 1'h0;
      write_enable_data_log_force[ 181] <= 1'h0;
      write_enable_data_log_force[ 182] <= 1'h0;
      write_enable_data_log_force[ 183] <= 1'h0;
      write_enable_data_log_force[ 184] <= 1'h0;
      write_enable_data_log_force[ 185] <= 1'h0;
      write_enable_data_log_force[ 186] <= 1'h0;
      write_enable_data_log_force[ 187] <= 1'h0;
      write_enable_data_log_force[ 188] <= 1'h0;
      write_enable_data_log_force[ 189] <= 1'h0;
      write_enable_data_log_force[ 190] <= 1'h0;
      write_enable_data_log_force[ 191] <= 1'h0;
      write_enable_data_log_force[ 192] <= 1'h0;
      write_enable_data_log_force[ 193] <= 1'h0;
      write_enable_data_log_force[ 194] <= 1'h0;
      write_enable_data_log_force[ 195] <= 1'h0;
      write_enable_data_log_force[ 196] <= 1'h0;
      write_enable_data_log_force[ 197] <= 1'h0;
      write_enable_data_log_force[ 198] <= 1'h0;
      write_enable_data_log_force[ 199] <= 1'h0;
      write_enable_data_log_force[ 200] <= 1'h0;
      write_enable_data_log_force[ 201] <= 1'h0;
      write_enable_data_log_force[ 202] <= 1'h0;
      write_enable_data_log_force[ 203] <= 1'h0;
      write_enable_data_log_force[ 204] <= 1'h0;
      write_enable_data_log_force[ 205] <= 1'h0;
      write_enable_data_log_force[ 206] <= 1'h0;
      write_enable_data_log_force[ 207] <= 1'h0;
      write_enable_data_log_force[ 208] <= 1'h0;
      write_enable_data_log_force[ 209] <= 1'h0;
      write_enable_data_log_force[ 210] <= 1'h0;
      write_enable_data_log_force[ 211] <= 1'h0;
      write_enable_data_log_force[ 212] <= 1'h0;
      write_enable_data_log_force[ 213] <= 1'h0;
      write_enable_data_log_force[ 214] <= 1'h0;
      write_enable_data_log_force[ 215] <= 1'h0;
      write_enable_data_log_force[ 216] <= 1'h0;
      write_enable_data_log_force[ 217] <= 1'h0;
      write_enable_data_log_force[ 218] <= 1'h0;
      write_enable_data_log_force[ 219] <= 1'h0;
      write_enable_data_log_force[ 220] <= 1'h0;
      write_enable_data_log_force[ 221] <= 1'h0;
      write_enable_data_log_force[ 222] <= 1'h0;
      write_enable_data_log_force[ 223] <= 1'h0;
      write_enable_data_log_force[ 224] <= 1'h0;
      write_enable_data_log_force[ 225] <= 1'h0;
      write_enable_data_log_force[ 226] <= 1'h0;
      write_enable_data_log_force[ 227] <= 1'h0;
      write_enable_data_log_force[ 228] <= 1'h0;
      write_enable_data_log_force[ 229] <= 1'h0;
      write_enable_data_log_force[ 230] <= 1'h0;
      write_enable_data_log_force[ 231] <= 1'h0;
      write_enable_data_log_force[ 232] <= 1'h0;
      write_enable_data_log_force[ 233] <= 1'h0;
      write_enable_data_log_force[ 234] <= 1'h0;
      write_enable_data_log_force[ 235] <= 1'h0;
      write_enable_data_log_force[ 236] <= 1'h0;
      write_enable_data_log_force[ 237] <= 1'h0;
      write_enable_data_log_force[ 238] <= 1'h0;
      write_enable_data_log_force[ 239] <= 1'h0;
      write_enable_data_log_force[ 240] <= 1'h0;
      write_enable_data_log_force[ 241] <= 1'h0;
      write_enable_data_log_force[ 242] <= 1'h0;
      write_enable_data_log_force[ 243] <= 1'h0;
      write_enable_data_log_force[ 244] <= 1'h0;
      write_enable_data_log_force[ 245] <= 1'h0;
      write_enable_data_log_force[ 246] <= 1'h0;
      write_enable_data_log_force[ 247] <= 1'h0;
      write_enable_data_log_force[ 248] <= 1'h0;
      write_enable_data_log_force[ 249] <= 1'h0;
      write_enable_data_log_force[ 250] <= 1'h0;
      write_enable_data_log_force[ 251] <= 1'h0;
      write_enable_data_log_force[ 252] <= 1'h0;
      write_enable_data_log_force[ 253] <= 1'h0;
      write_enable_data_log_force[ 254] <= 1'h0;
      write_enable_data_log_force[ 255] <= 1'h0;
      write_enable_data_log_force[ 256] <= 1'h0;
      write_enable_data_log_force[ 257] <= 1'h0;
      write_enable_data_log_force[ 258] <= 1'h0;
      write_enable_data_log_force[ 259] <= 1'h0;
      write_enable_data_log_force[ 260] <= 1'h0;
      write_enable_data_log_force[ 261] <= 1'h0;
      write_enable_data_log_force[ 262] <= 1'h0;
      write_enable_data_log_force[ 263] <= 1'h0;
      write_enable_data_log_force[ 264] <= 1'h0;
      write_enable_data_log_force[ 265] <= 1'h0;
      write_enable_data_log_force[ 266] <= 1'h0;
      write_enable_data_log_force[ 267] <= 1'h0;
      write_enable_data_log_force[ 268] <= 1'h0;
      write_enable_data_log_force[ 269] <= 1'h0;
      write_enable_data_log_force[ 270] <= 1'h0;
      write_enable_data_log_force[ 271] <= 1'h0;
      write_enable_data_log_force[ 272] <= 1'h0;
      write_enable_data_log_force[ 273] <= 1'h0;
      write_enable_data_log_force[ 274] <= 1'h0;
      write_enable_data_log_force[ 275] <= 1'h0;
      write_enable_data_log_force[ 276] <= 1'h0;
      write_enable_data_log_force[ 277] <= 1'h0;
      write_enable_data_log_force[ 278] <= 1'h0;
      write_enable_data_log_force[ 279] <= 1'h0;
      write_enable_data_log_force[ 280] <= 1'h0;
      write_enable_data_log_force[ 281] <= 1'h0;
      write_enable_data_log_force[ 282] <= 1'h0;
      write_enable_data_log_force[ 283] <= 1'h0;
      write_enable_data_log_force[ 284] <= 1'h0;
      write_enable_data_log_force[ 285] <= 1'h0;
      write_enable_data_log_force[ 286] <= 1'h0;
      write_enable_data_log_force[ 287] <= 1'h0;
      write_enable_data_log_force[ 288] <= 1'h0;
      write_enable_data_log_force[ 289] <= 1'h0;
      write_enable_data_log_force[ 290] <= 1'h0;
      write_enable_data_log_force[ 291] <= 1'h0;
      write_enable_data_log_force[ 292] <= 1'h0;
      write_enable_data_log_force[ 293] <= 1'h0;
      write_enable_data_log_force[ 294] <= 1'h0;
      write_enable_data_log_force[ 295] <= 1'h0;
      write_enable_data_log_force[ 296] <= 1'h0;
      write_enable_data_log_force[ 297] <= 1'h0;
      write_enable_data_log_force[ 298] <= 1'h0;
      write_enable_data_log_force[ 299] <= 1'h0;
      write_enable_data_log_force[ 300] <= 1'h0;
      write_enable_data_log_force[ 301] <= 1'h0;
      write_enable_data_log_force[ 302] <= 1'h0;
      write_enable_data_log_force[ 303] <= 1'h0;
      write_enable_data_log_force[ 304] <= 1'h0;
      write_enable_data_log_force[ 305] <= 1'h0;
      write_enable_data_log_force[ 306] <= 1'h0;
      write_enable_data_log_force[ 307] <= 1'h0;
      write_enable_data_log_force[ 308] <= 1'h0;
      write_enable_data_log_force[ 309] <= 1'h0;
      write_enable_data_log_force[ 310] <= 1'h0;
      write_enable_data_log_force[ 311] <= 1'h0;
      write_enable_data_log_force[ 312] <= 1'h0;
      write_enable_data_log_force[ 313] <= 1'h0;
      write_enable_data_log_force[ 314] <= 1'h0;
      write_enable_data_log_force[ 315] <= 1'h0;
      write_enable_data_log_force[ 316] <= 1'h0;
      write_enable_data_log_force[ 317] <= 1'h0;
      write_enable_data_log_force[ 318] <= 1'h0;
      write_enable_data_log_force[ 319] <= 1'h0;
      write_enable_data_log_force[ 320] <= 1'h0;
      write_enable_data_log_force[ 321] <= 1'h0;
      write_enable_data_log_force[ 322] <= 1'h0;
      write_enable_data_log_force[ 323] <= 1'h0;
      write_enable_data_log_force[ 324] <= 1'h0;
      write_enable_data_log_force[ 325] <= 1'h0;
      write_enable_data_log_force[ 326] <= 1'h0;
      write_enable_data_log_force[ 327] <= 1'h0;
      write_enable_data_log_force[ 328] <= 1'h0;
      write_enable_data_log_force[ 329] <= 1'h0;
      write_enable_data_log_force[ 330] <= 1'h0;
      write_enable_data_log_force[ 331] <= 1'h0;
      write_enable_data_log_force[ 332] <= 1'h0;
      write_enable_data_log_force[ 333] <= 1'h0;
      write_enable_data_log_force[ 334] <= 1'h0;
      write_enable_data_log_force[ 335] <= 1'h0;
      write_enable_data_log_force[ 336] <= 1'h0;
      write_enable_data_log_force[ 337] <= 1'h0;
      write_enable_data_log_force[ 338] <= 1'h0;
      write_enable_data_log_force[ 339] <= 1'h0;
      write_enable_data_log_force[ 340] <= 1'h0;
      write_enable_data_log_force[ 341] <= 1'h0;
      write_enable_data_log_force[ 342] <= 1'h0;
      write_enable_data_log_force[ 343] <= 1'h0;
      write_enable_data_log_force[ 344] <= 1'h0;
      write_enable_data_log_force[ 345] <= 1'h0;
      write_enable_data_log_force[ 346] <= 1'h0;
      write_enable_data_log_force[ 347] <= 1'h0;
      write_enable_data_log_force[ 348] <= 1'h0;
      write_enable_data_log_force[ 349] <= 1'h0;
      write_enable_data_log_force[ 350] <= 1'h0;
      write_enable_data_log_force[ 351] <= 1'h0;
      write_enable_data_log_force[ 352] <= 1'h0;
      write_enable_data_log_force[ 353] <= 1'h0;
      write_enable_data_log_force[ 354] <= 1'h0;
      write_enable_data_log_force[ 355] <= 1'h0;
      write_enable_data_log_force[ 356] <= 1'h0;
      write_enable_data_log_force[ 357] <= 1'h0;
      write_enable_data_log_force[ 358] <= 1'h0;
      write_enable_data_log_force[ 359] <= 1'h0;
      write_enable_data_log_force[ 360] <= 1'h0;
      write_enable_data_log_force[ 361] <= 1'h0;
      write_enable_data_log_force[ 362] <= 1'h0;
      write_enable_data_log_force[ 363] <= 1'h0;
      write_enable_data_log_force[ 364] <= 1'h0;
      write_enable_data_log_force[ 365] <= 1'h0;
      write_enable_data_log_force[ 366] <= 1'h0;
      write_enable_data_log_force[ 367] <= 1'h0;
      write_enable_data_log_force[ 368] <= 1'h0;
      write_enable_data_log_force[ 369] <= 1'h0;
      write_enable_data_log_force[ 370] <= 1'h0;
      write_enable_data_log_force[ 371] <= 1'h0;
      write_enable_data_log_force[ 372] <= 1'h0;
      write_enable_data_log_force[ 373] <= 1'h0;
      write_enable_data_log_force[ 374] <= 1'h0;
      write_enable_data_log_force[ 375] <= 1'h0;
      write_enable_data_log_force[ 376] <= 1'h0;
      write_enable_data_log_force[ 377] <= 1'h0;
      write_enable_data_log_force[ 378] <= 1'h0;
      write_enable_data_log_force[ 379] <= 1'h0;
      write_enable_data_log_force[ 380] <= 1'h0;
      write_enable_data_log_force[ 381] <= 1'h0;
      write_enable_data_log_force[ 382] <= 1'h0;
      write_enable_data_log_force[ 383] <= 1'h0;
      write_enable_data_log_force[ 384] <= 1'h0;
      write_enable_data_log_force[ 385] <= 1'h0;
      write_enable_data_log_force[ 386] <= 1'h0;
      write_enable_data_log_force[ 387] <= 1'h0;
      write_enable_data_log_force[ 388] <= 1'h0;
      write_enable_data_log_force[ 389] <= 1'h0;
      write_enable_data_log_force[ 390] <= 1'h0;
      write_enable_data_log_force[ 391] <= 1'h0;
      write_enable_data_log_force[ 392] <= 1'h0;
      write_enable_data_log_force[ 393] <= 1'h0;
      write_enable_data_log_force[ 394] <= 1'h0;
      write_enable_data_log_force[ 395] <= 1'h0;
      write_enable_data_log_force[ 396] <= 1'h0;
      write_enable_data_log_force[ 397] <= 1'h0;
      write_enable_data_log_force[ 398] <= 1'h0;
      write_enable_data_log_force[ 399] <= 1'h0;
      write_enable_data_log_force[ 400] <= 1'h0;
      write_enable_data_log_force[ 401] <= 1'h0;
      write_enable_data_log_force[ 402] <= 1'h0;
      write_enable_data_log_force[ 403] <= 1'h0;
      write_enable_data_log_force[ 404] <= 1'h0;
      write_enable_data_log_force[ 405] <= 1'h0;
      write_enable_data_log_force[ 406] <= 1'h0;
      write_enable_data_log_force[ 407] <= 1'h0;
      write_enable_data_log_force[ 408] <= 1'h0;
      write_enable_data_log_force[ 409] <= 1'h0;
      write_enable_data_log_force[ 410] <= 1'h0;
      write_enable_data_log_force[ 411] <= 1'h0;
      write_enable_data_log_force[ 412] <= 1'h0;
      write_enable_data_log_force[ 413] <= 1'h0;
      write_enable_data_log_force[ 414] <= 1'h0;
      write_enable_data_log_force[ 415] <= 1'h0;
      write_enable_data_log_force[ 416] <= 1'h0;
      write_enable_data_log_force[ 417] <= 1'h0;
      write_enable_data_log_force[ 418] <= 1'h0;
      write_enable_data_log_force[ 419] <= 1'h0;
      write_enable_data_log_force[ 420] <= 1'h0;
      write_enable_data_log_force[ 421] <= 1'h0;
      write_enable_data_log_force[ 422] <= 1'h0;
      write_enable_data_log_force[ 423] <= 1'h0;
      write_enable_data_log_force[ 424] <= 1'h0;
      write_enable_data_log_force[ 425] <= 1'h0;
      write_enable_data_log_force[ 426] <= 1'h0;
      write_enable_data_log_force[ 427] <= 1'h0;
      write_enable_data_log_force[ 428] <= 1'h0;
      write_enable_data_log_force[ 429] <= 1'h0;
      write_enable_data_log_force[ 430] <= 1'h0;
      write_enable_data_log_force[ 431] <= 1'h0;
      write_enable_data_log_force[ 432] <= 1'h0;
      write_enable_data_log_force[ 433] <= 1'h0;
      write_enable_data_log_force[ 434] <= 1'h0;
      write_enable_data_log_force[ 435] <= 1'h0;
      write_enable_data_log_force[ 436] <= 1'h0;
      write_enable_data_log_force[ 437] <= 1'h0;
      write_enable_data_log_force[ 438] <= 1'h0;
      write_enable_data_log_force[ 439] <= 1'h0;
      write_enable_data_log_force[ 440] <= 1'h0;
      write_enable_data_log_force[ 441] <= 1'h0;
      write_enable_data_log_force[ 442] <= 1'h0;
      write_enable_data_log_force[ 443] <= 1'h0;
      write_enable_data_log_force[ 444] <= 1'h0;
      write_enable_data_log_force[ 445] <= 1'h0;
      write_enable_data_log_force[ 446] <= 1'h0;
      write_enable_data_log_force[ 447] <= 1'h0;
      write_enable_data_log_force[ 448] <= 1'h0;
      write_enable_data_log_force[ 449] <= 1'h0;
      write_enable_data_log_force[ 450] <= 1'h0;
      write_enable_data_log_force[ 451] <= 1'h0;
      write_enable_data_log_force[ 452] <= 1'h0;
      write_enable_data_log_force[ 453] <= 1'h0;
      write_enable_data_log_force[ 454] <= 1'h0;
      write_enable_data_log_force[ 455] <= 1'h0;
      write_enable_data_log_force[ 456] <= 1'h0;
      write_enable_data_log_force[ 457] <= 1'h0;
      write_enable_data_log_force[ 458] <= 1'h0;
      write_enable_data_log_force[ 459] <= 1'h0;
      write_enable_data_log_force[ 460] <= 1'h0;
      write_enable_data_log_force[ 461] <= 1'h0;
      write_enable_data_log_force[ 462] <= 1'h0;
      write_enable_data_log_force[ 463] <= 1'h0;
      write_enable_data_log_force[ 464] <= 1'h0;
      write_enable_data_log_force[ 465] <= 1'h0;
      write_enable_data_log_force[ 466] <= 1'h0;
      write_enable_data_log_force[ 467] <= 1'h0;
      write_enable_data_log_force[ 468] <= 1'h0;
      write_enable_data_log_force[ 469] <= 1'h0;
      write_enable_data_log_force[ 470] <= 1'h0;
      write_enable_data_log_force[ 471] <= 1'h0;
      write_enable_data_log_force[ 472] <= 1'h0;
      write_enable_data_log_force[ 473] <= 1'h0;
      write_enable_data_log_force[ 474] <= 1'h0;
      write_enable_data_log_force[ 475] <= 1'h0;
      write_enable_data_log_force[ 476] <= 1'h0;
      write_enable_data_log_force[ 477] <= 1'h0;
      write_enable_data_log_force[ 478] <= 1'h0;
      write_enable_data_log_force[ 479] <= 1'h0;
      write_enable_data_log_force[ 480] <= 1'h0;
      write_enable_data_log_force[ 481] <= 1'h0;
      write_enable_data_log_force[ 482] <= 1'h0;
      write_enable_data_log_force[ 483] <= 1'h0;
      write_enable_data_log_force[ 484] <= 1'h0;
      write_enable_data_log_force[ 485] <= 1'h0;
      write_enable_data_log_force[ 486] <= 1'h0;
      write_enable_data_log_force[ 487] <= 1'h0;
      write_enable_data_log_force[ 488] <= 1'h0;
      write_enable_data_log_force[ 489] <= 1'h0;
      write_enable_data_log_force[ 490] <= 1'h0;
      write_enable_data_log_force[ 491] <= 1'h0;
      write_enable_data_log_force[ 492] <= 1'h0;
      write_enable_data_log_force[ 493] <= 1'h0;
      write_enable_data_log_force[ 494] <= 1'h0;
      write_enable_data_log_force[ 495] <= 1'h0;
      write_enable_data_log_force[ 496] <= 1'h0;
      write_enable_data_log_force[ 497] <= 1'h0;
      write_enable_data_log_force[ 498] <= 1'h0;
      write_enable_data_log_force[ 499] <= 1'h0;
      write_enable_data_log_force[ 500] <= 1'h0;
      write_enable_data_log_force[ 501] <= 1'h0;
      write_enable_data_log_force[ 502] <= 1'h0;
      write_enable_data_log_force[ 503] <= 1'h0;
      write_enable_data_log_force[ 504] <= 1'h0;
      write_enable_data_log_force[ 505] <= 1'h0;
      write_enable_data_log_force[ 506] <= 1'h0;
      write_enable_data_log_force[ 507] <= 1'h0;
      write_enable_data_log_force[ 508] <= 1'h0;
      write_enable_data_log_force[ 509] <= 1'h0;
      write_enable_data_log_force[ 510] <= 1'h0;
      write_enable_data_log_force[ 511] <= 1'h0;
      write_enable_data_log_force[ 512] <= 1'h0;
      write_enable_data_log_force[ 513] <= 1'h0;
      write_enable_data_log_force[ 514] <= 1'h0;
      write_enable_data_log_force[ 515] <= 1'h0;
      write_enable_data_log_force[ 516] <= 1'h0;
      write_enable_data_log_force[ 517] <= 1'h0;
      write_enable_data_log_force[ 518] <= 1'h0;
      write_enable_data_log_force[ 519] <= 1'h0;
      write_enable_data_log_force[ 520] <= 1'h0;
      write_enable_data_log_force[ 521] <= 1'h0;
      write_enable_data_log_force[ 522] <= 1'h0;
      write_enable_data_log_force[ 523] <= 1'h0;
      write_enable_data_log_force[ 524] <= 1'h0;
      write_enable_data_log_force[ 525] <= 1'h0;
      write_enable_data_log_force[ 526] <= 1'h0;
      write_enable_data_log_force[ 527] <= 1'h0;
      write_enable_data_log_force[ 528] <= 1'h0;
      write_enable_data_log_force[ 529] <= 1'h0;
      write_enable_data_log_force[ 530] <= 1'h0;
      write_enable_data_log_force[ 531] <= 1'h0;
      write_enable_data_log_force[ 532] <= 1'h0;
      write_enable_data_log_force[ 533] <= 1'h0;
      write_enable_data_log_force[ 534] <= 1'h0;
      write_enable_data_log_force[ 535] <= 1'h0;
      write_enable_data_log_force[ 536] <= 1'h0;
      write_enable_data_log_force[ 537] <= 1'h0;
      write_enable_data_log_force[ 538] <= 1'h0;
      write_enable_data_log_force[ 539] <= 1'h0;
      write_enable_data_log_force[ 540] <= 1'h0;
      write_enable_data_log_force[ 541] <= 1'h0;
      write_enable_data_log_force[ 542] <= 1'h0;
      write_enable_data_log_force[ 543] <= 1'h0;
      write_enable_data_log_force[ 544] <= 1'h0;
      write_enable_data_log_force[ 545] <= 1'h0;
      write_enable_data_log_force[ 546] <= 1'h0;
      write_enable_data_log_force[ 547] <= 1'h0;
      write_enable_data_log_force[ 548] <= 1'h0;
      write_enable_data_log_force[ 549] <= 1'h0;
      write_enable_data_log_force[ 550] <= 1'h0;
      write_enable_data_log_force[ 551] <= 1'h0;
      write_enable_data_log_force[ 552] <= 1'h0;
      write_enable_data_log_force[ 553] <= 1'h0;
      write_enable_data_log_force[ 554] <= 1'h0;
      write_enable_data_log_force[ 555] <= 1'h0;
      write_enable_data_log_force[ 556] <= 1'h0;
      write_enable_data_log_force[ 557] <= 1'h0;
      write_enable_data_log_force[ 558] <= 1'h0;
      write_enable_data_log_force[ 559] <= 1'h0;
      write_enable_data_log_force[ 560] <= 1'h0;
      write_enable_data_log_force[ 561] <= 1'h0;
      write_enable_data_log_force[ 562] <= 1'h0;
      write_enable_data_log_force[ 563] <= 1'h0;
      write_enable_data_log_force[ 564] <= 1'h0;
      write_enable_data_log_force[ 565] <= 1'h0;
      write_enable_data_log_force[ 566] <= 1'h0;
      write_enable_data_log_force[ 567] <= 1'h0;
      write_enable_data_log_force[ 568] <= 1'h0;
      write_enable_data_log_force[ 569] <= 1'h0;
      write_enable_data_log_force[ 570] <= 1'h0;
      write_enable_data_log_force[ 571] <= 1'h0;
      write_enable_data_log_force[ 572] <= 1'h0;
      write_enable_data_log_force[ 573] <= 1'h0;
      write_enable_data_log_force[ 574] <= 1'h0;
      write_enable_data_log_force[ 575] <= 1'h0;
      write_enable_data_log_force[ 576] <= 1'h0;
      write_enable_data_log_force[ 577] <= 1'h0;
      write_enable_data_log_force[ 578] <= 1'h0;
      write_enable_data_log_force[ 579] <= 1'h0;
      write_enable_data_log_force[ 580] <= 1'h0;
      write_enable_data_log_force[ 581] <= 1'h0;
      write_enable_data_log_force[ 582] <= 1'h0;
      write_enable_data_log_force[ 583] <= 1'h0;
      write_enable_data_log_force[ 584] <= 1'h0;
      write_enable_data_log_force[ 585] <= 1'h0;
      write_enable_data_log_force[ 586] <= 1'h0;
      write_enable_data_log_force[ 587] <= 1'h0;
      write_enable_data_log_force[ 588] <= 1'h0;
      write_enable_data_log_force[ 589] <= 1'h0;
      write_enable_data_log_force[ 590] <= 1'h0;
      write_enable_data_log_force[ 591] <= 1'h0;
      write_enable_data_log_force[ 592] <= 1'h0;
      write_enable_data_log_force[ 593] <= 1'h0;
      write_enable_data_log_force[ 594] <= 1'h0;
      write_enable_data_log_force[ 595] <= 1'h0;
      write_enable_data_log_force[ 596] <= 1'h0;
      write_enable_data_log_force[ 597] <= 1'h0;
      write_enable_data_log_force[ 598] <= 1'h0;
      write_enable_data_log_force[ 599] <= 1'h0;
      write_enable_data_log_force[ 600] <= 1'h0;
      write_enable_data_log_force[ 601] <= 1'h0;
      write_enable_data_log_force[ 602] <= 1'h0;
      write_enable_data_log_force[ 603] <= 1'h0;
      write_enable_data_log_force[ 604] <= 1'h0;
      write_enable_data_log_force[ 605] <= 1'h0;
      write_enable_data_log_force[ 606] <= 1'h0;
      write_enable_data_log_force[ 607] <= 1'h0;
      write_enable_data_log_force[ 608] <= 1'h0;
      write_enable_data_log_force[ 609] <= 1'h0;
      write_enable_data_log_force[ 610] <= 1'h0;
      write_enable_data_log_force[ 611] <= 1'h0;
      write_enable_data_log_force[ 612] <= 1'h0;
      write_enable_data_log_force[ 613] <= 1'h0;
      write_enable_data_log_force[ 614] <= 1'h0;
      write_enable_data_log_force[ 615] <= 1'h0;
      write_enable_data_log_force[ 616] <= 1'h0;
      write_enable_data_log_force[ 617] <= 1'h0;
      write_enable_data_log_force[ 618] <= 1'h0;
      write_enable_data_log_force[ 619] <= 1'h0;
      write_enable_data_log_force[ 620] <= 1'h0;
      write_enable_data_log_force[ 621] <= 1'h0;
      write_enable_data_log_force[ 622] <= 1'h0;
      write_enable_data_log_force[ 623] <= 1'h0;
      write_enable_data_log_force[ 624] <= 1'h0;
      write_enable_data_log_force[ 625] <= 1'h0;
      write_enable_data_log_force[ 626] <= 1'h0;
      write_enable_data_log_force[ 627] <= 1'h0;
      write_enable_data_log_force[ 628] <= 1'h0;
      write_enable_data_log_force[ 629] <= 1'h0;
      write_enable_data_log_force[ 630] <= 1'h0;
      write_enable_data_log_force[ 631] <= 1'h0;
      write_enable_data_log_force[ 632] <= 1'h0;
      write_enable_data_log_force[ 633] <= 1'h0;
      write_enable_data_log_force[ 634] <= 1'h0;
      write_enable_data_log_force[ 635] <= 1'h0;
      write_enable_data_log_force[ 636] <= 1'h0;
      write_enable_data_log_force[ 637] <= 1'h0;
      write_enable_data_log_force[ 638] <= 1'h0;
      write_enable_data_log_force[ 639] <= 1'h0;
      write_enable_data_log_force[ 640] <= 1'h0;
      write_enable_data_log_force[ 641] <= 1'h0;
      write_enable_data_log_force[ 642] <= 1'h0;
      write_enable_data_log_force[ 643] <= 1'h0;
      write_enable_data_log_force[ 644] <= 1'h0;
      write_enable_data_log_force[ 645] <= 1'h0;
      write_enable_data_log_force[ 646] <= 1'h0;
      write_enable_data_log_force[ 647] <= 1'h0;
      write_enable_data_log_force[ 648] <= 1'h0;
      write_enable_data_log_force[ 649] <= 1'h0;
      write_enable_data_log_force[ 650] <= 1'h0;
      write_enable_data_log_force[ 651] <= 1'h0;
      write_enable_data_log_force[ 652] <= 1'h0;
      write_enable_data_log_force[ 653] <= 1'h0;
      write_enable_data_log_force[ 654] <= 1'h0;
      write_enable_data_log_force[ 655] <= 1'h0;
      write_enable_data_log_force[ 656] <= 1'h0;
      write_enable_data_log_force[ 657] <= 1'h0;
      write_enable_data_log_force[ 658] <= 1'h0;
      write_enable_data_log_force[ 659] <= 1'h0;
      write_enable_data_log_force[ 660] <= 1'h0;
      write_enable_data_log_force[ 661] <= 1'h0;
      write_enable_data_log_force[ 662] <= 1'h0;
      write_enable_data_log_force[ 663] <= 1'h0;
      write_enable_data_log_force[ 664] <= 1'h0;
      write_enable_data_log_force[ 665] <= 1'h0;
      write_enable_data_log_force[ 666] <= 1'h0;
      write_enable_data_log_force[ 667] <= 1'h0;
      write_enable_data_log_force[ 668] <= 1'h0;
      write_enable_data_log_force[ 669] <= 1'h0;
      write_enable_data_log_force[ 670] <= 1'h0;
      write_enable_data_log_force[ 671] <= 1'h0;
      write_enable_data_log_force[ 672] <= 1'h0;
      write_enable_data_log_force[ 673] <= 1'h0;
      write_enable_data_log_force[ 674] <= 1'h0;
      write_enable_data_log_force[ 675] <= 1'h0;
      write_enable_data_log_force[ 676] <= 1'h0;
      write_enable_data_log_force[ 677] <= 1'h0;
      write_enable_data_log_force[ 678] <= 1'h0;
      write_enable_data_log_force[ 679] <= 1'h0;
      write_enable_data_log_force[ 680] <= 1'h0;
      write_enable_data_log_force[ 681] <= 1'h0;
      write_enable_data_log_force[ 682] <= 1'h0;
      write_enable_data_log_force[ 683] <= 1'h0;
      write_enable_data_log_force[ 684] <= 1'h0;
      write_enable_data_log_force[ 685] <= 1'h0;
      write_enable_data_log_force[ 686] <= 1'h0;
      write_enable_data_log_force[ 687] <= 1'h0;
      write_enable_data_log_force[ 688] <= 1'h0;
      write_enable_data_log_force[ 689] <= 1'h0;
      write_enable_data_log_force[ 690] <= 1'h0;
      write_enable_data_log_force[ 691] <= 1'h0;
      write_enable_data_log_force[ 692] <= 1'h0;
      write_enable_data_log_force[ 693] <= 1'h0;
      write_enable_data_log_force[ 694] <= 1'h0;
      write_enable_data_log_force[ 695] <= 1'h0;
      write_enable_data_log_force[ 696] <= 1'h0;
      write_enable_data_log_force[ 697] <= 1'h0;
      write_enable_data_log_force[ 698] <= 1'h0;
      write_enable_data_log_force[ 699] <= 1'h0;
      write_enable_data_log_force[ 700] <= 1'h0;
      write_enable_data_log_force[ 701] <= 1'h0;
      write_enable_data_log_force[ 702] <= 1'h0;
      write_enable_data_log_force[ 703] <= 1'h0;
      write_enable_data_log_force[ 704] <= 1'h0;
      write_enable_data_log_force[ 705] <= 1'h0;
      write_enable_data_log_force[ 706] <= 1'h0;
      write_enable_data_log_force[ 707] <= 1'h0;
      write_enable_data_log_force[ 708] <= 1'h0;
      write_enable_data_log_force[ 709] <= 1'h0;
      write_enable_data_log_force[ 710] <= 1'h0;
      write_enable_data_log_force[ 711] <= 1'h0;
      write_enable_data_log_force[ 712] <= 1'h0;
      write_enable_data_log_force[ 713] <= 1'h0;
      write_enable_data_log_force[ 714] <= 1'h0;
      write_enable_data_log_force[ 715] <= 1'h0;
      write_enable_data_log_force[ 716] <= 1'h0;
      write_enable_data_log_force[ 717] <= 1'h0;
      write_enable_data_log_force[ 718] <= 1'h0;
      write_enable_data_log_force[ 719] <= 1'h0;
      write_enable_data_log_force[ 720] <= 1'h0;
      write_enable_data_log_force[ 721] <= 1'h0;
      write_enable_data_log_force[ 722] <= 1'h0;
      write_enable_data_log_force[ 723] <= 1'h0;
      write_enable_data_log_force[ 724] <= 1'h0;
      write_enable_data_log_force[ 725] <= 1'h0;
      write_enable_data_log_force[ 726] <= 1'h0;
      write_enable_data_log_force[ 727] <= 1'h0;
      write_enable_data_log_force[ 728] <= 1'h0;
      write_enable_data_log_force[ 729] <= 1'h0;
      write_enable_data_log_force[ 730] <= 1'h0;
      write_enable_data_log_force[ 731] <= 1'h0;
      write_enable_data_log_force[ 732] <= 1'h0;
      write_enable_data_log_force[ 733] <= 1'h0;
      write_enable_data_log_force[ 734] <= 1'h0;
      write_enable_data_log_force[ 735] <= 1'h0;
      write_enable_data_log_force[ 736] <= 1'h0;
      write_enable_data_log_force[ 737] <= 1'h0;
      write_enable_data_log_force[ 738] <= 1'h0;
      write_enable_data_log_force[ 739] <= 1'h0;
      write_enable_data_log_force[ 740] <= 1'h0;
      write_enable_data_log_force[ 741] <= 1'h0;
      write_enable_data_log_force[ 742] <= 1'h0;
      write_enable_data_log_force[ 743] <= 1'h0;
      write_enable_data_log_force[ 744] <= 1'h0;
      write_enable_data_log_force[ 745] <= 1'h0;
      write_enable_data_log_force[ 746] <= 1'h0;
      write_enable_data_log_force[ 747] <= 1'h0;
      write_enable_data_log_force[ 748] <= 1'h0;
      write_enable_data_log_force[ 749] <= 1'h0;
      write_enable_data_log_force[ 750] <= 1'h0;
      write_enable_data_log_force[ 751] <= 1'h0;
      write_enable_data_log_force[ 752] <= 1'h0;
      write_enable_data_log_force[ 753] <= 1'h0;
      write_enable_data_log_force[ 754] <= 1'h0;
      write_enable_data_log_force[ 755] <= 1'h0;
      write_enable_data_log_force[ 756] <= 1'h0;
      write_enable_data_log_force[ 757] <= 1'h0;
      write_enable_data_log_force[ 758] <= 1'h0;
      write_enable_data_log_force[ 759] <= 1'h0;
      write_enable_data_log_force[ 760] <= 1'h0;
      write_enable_data_log_force[ 761] <= 1'h0;
      write_enable_data_log_force[ 762] <= 1'h0;
      write_enable_data_log_force[ 763] <= 1'h0;
      write_enable_data_log_force[ 764] <= 1'h0;
      write_enable_data_log_force[ 765] <= 1'h0;
      write_enable_data_log_force[ 766] <= 1'h0;
      write_enable_data_log_force[ 767] <= 1'h0;
      write_enable_data_log_force[ 768] <= 1'h0;
      write_enable_data_log_force[ 769] <= 1'h0;
      write_enable_data_log_force[ 770] <= 1'h0;
      write_enable_data_log_force[ 771] <= 1'h0;
      write_enable_data_log_force[ 772] <= 1'h0;
      write_enable_data_log_force[ 773] <= 1'h0;
      write_enable_data_log_force[ 774] <= 1'h0;
      write_enable_data_log_force[ 775] <= 1'h0;
      write_enable_data_log_force[ 776] <= 1'h0;
      write_enable_data_log_force[ 777] <= 1'h0;
      write_enable_data_log_force[ 778] <= 1'h0;
      write_enable_data_log_force[ 779] <= 1'h0;
      write_enable_data_log_force[ 780] <= 1'h0;
      write_enable_data_log_force[ 781] <= 1'h0;
      write_enable_data_log_force[ 782] <= 1'h0;
      write_enable_data_log_force[ 783] <= 1'h0;
      write_enable_data_log_force[ 784] <= 1'h0;
      write_enable_data_log_force[ 785] <= 1'h0;
      write_enable_data_log_force[ 786] <= 1'h0;
      write_enable_data_log_force[ 787] <= 1'h0;
      write_enable_data_log_force[ 788] <= 1'h0;
      write_enable_data_log_force[ 789] <= 1'h0;
      write_enable_data_log_force[ 790] <= 1'h0;
      write_enable_data_log_force[ 791] <= 1'h0;
      write_enable_data_log_force[ 792] <= 1'h0;
      write_enable_data_log_force[ 793] <= 1'h0;
      write_enable_data_log_force[ 794] <= 1'h0;
      write_enable_data_log_force[ 795] <= 1'h0;
      write_enable_data_log_force[ 796] <= 1'h0;
      write_enable_data_log_force[ 797] <= 1'h0;
      write_enable_data_log_force[ 798] <= 1'h0;
      write_enable_data_log_force[ 799] <= 1'h0;
      write_enable_data_log_force[ 800] <= 1'h0;
      write_enable_data_log_force[ 801] <= 1'h0;
      write_enable_data_log_force[ 802] <= 1'h0;
      write_enable_data_log_force[ 803] <= 1'h0;
      write_enable_data_log_force[ 804] <= 1'h0;
      write_enable_data_log_force[ 805] <= 1'h0;
      write_enable_data_log_force[ 806] <= 1'h0;
      write_enable_data_log_force[ 807] <= 1'h0;
      write_enable_data_log_force[ 808] <= 1'h0;
      write_enable_data_log_force[ 809] <= 1'h0;
      write_enable_data_log_force[ 810] <= 1'h0;
      write_enable_data_log_force[ 811] <= 1'h0;
      write_enable_data_log_force[ 812] <= 1'h0;
      write_enable_data_log_force[ 813] <= 1'h0;
      write_enable_data_log_force[ 814] <= 1'h0;
      write_enable_data_log_force[ 815] <= 1'h0;
      write_enable_data_log_force[ 816] <= 1'h0;
      write_enable_data_log_force[ 817] <= 1'h0;
      write_enable_data_log_force[ 818] <= 1'h0;
      write_enable_data_log_force[ 819] <= 1'h0;
      write_enable_data_log_force[ 820] <= 1'h0;
      write_enable_data_log_force[ 821] <= 1'h0;
      write_enable_data_log_force[ 822] <= 1'h0;
      write_enable_data_log_force[ 823] <= 1'h0;
      write_enable_data_log_force[ 824] <= 1'h0;
      write_enable_data_log_force[ 825] <= 1'h0;
      write_enable_data_log_force[ 826] <= 1'h0;
      write_enable_data_log_force[ 827] <= 1'h0;
      write_enable_data_log_force[ 828] <= 1'h0;
      write_enable_data_log_force[ 829] <= 1'h0;
      write_enable_data_log_force[ 830] <= 1'h0;
      write_enable_data_log_force[ 831] <= 1'h0;
      write_enable_data_log_force[ 832] <= 1'h0;
      write_enable_data_log_force[ 833] <= 1'h0;
      write_enable_data_log_force[ 834] <= 1'h0;
      write_enable_data_log_force[ 835] <= 1'h0;
      write_enable_data_log_force[ 836] <= 1'h0;
      write_enable_data_log_force[ 837] <= 1'h0;
      write_enable_data_log_force[ 838] <= 1'h0;
      write_enable_data_log_force[ 839] <= 1'h0;
      write_enable_data_log_force[ 840] <= 1'h0;
      write_enable_data_log_force[ 841] <= 1'h0;
      write_enable_data_log_force[ 842] <= 1'h0;
      write_enable_data_log_force[ 843] <= 1'h0;
      write_enable_data_log_force[ 844] <= 1'h0;
      write_enable_data_log_force[ 845] <= 1'h0;
      write_enable_data_log_force[ 846] <= 1'h0;
      write_enable_data_log_force[ 847] <= 1'h0;
      write_enable_data_log_force[ 848] <= 1'h0;
      write_enable_data_log_force[ 849] <= 1'h0;
      write_enable_data_log_force[ 850] <= 1'h0;
      write_enable_data_log_force[ 851] <= 1'h0;
      write_enable_data_log_force[ 852] <= 1'h0;
      write_enable_data_log_force[ 853] <= 1'h0;
      write_enable_data_log_force[ 854] <= 1'h0;
      write_enable_data_log_force[ 855] <= 1'h0;
      write_enable_data_log_force[ 856] <= 1'h0;
      write_enable_data_log_force[ 857] <= 1'h0;
      write_enable_data_log_force[ 858] <= 1'h0;
      write_enable_data_log_force[ 859] <= 1'h0;
      write_enable_data_log_force[ 860] <= 1'h0;
      write_enable_data_log_force[ 861] <= 1'h0;
      write_enable_data_log_force[ 862] <= 1'h0;
      write_enable_data_log_force[ 863] <= 1'h0;
      write_enable_data_log_force[ 864] <= 1'h0;
      write_enable_data_log_force[ 865] <= 1'h0;
      write_enable_data_log_force[ 866] <= 1'h0;
      write_enable_data_log_force[ 867] <= 1'h0;
      write_enable_data_log_force[ 868] <= 1'h0;
      write_enable_data_log_force[ 869] <= 1'h0;
      write_enable_data_log_force[ 870] <= 1'h0;
      write_enable_data_log_force[ 871] <= 1'h0;
      write_enable_data_log_force[ 872] <= 1'h0;
      write_enable_data_log_force[ 873] <= 1'h0;
      write_enable_data_log_force[ 874] <= 1'h0;
      write_enable_data_log_force[ 875] <= 1'h0;
      write_enable_data_log_force[ 876] <= 1'h0;
      write_enable_data_log_force[ 877] <= 1'h0;
      write_enable_data_log_force[ 878] <= 1'h0;
      write_enable_data_log_force[ 879] <= 1'h0;
      write_enable_data_log_force[ 880] <= 1'h0;
      write_enable_data_log_force[ 881] <= 1'h0;
      write_enable_data_log_force[ 882] <= 1'h0;
      write_enable_data_log_force[ 883] <= 1'h0;
      write_enable_data_log_force[ 884] <= 1'h0;
      write_enable_data_log_force[ 885] <= 1'h0;
      write_enable_data_log_force[ 886] <= 1'h0;
      write_enable_data_log_force[ 887] <= 1'h0;
      write_enable_data_log_force[ 888] <= 1'h0;
      write_enable_data_log_force[ 889] <= 1'h0;
      write_enable_data_log_force[ 890] <= 1'h0;
      write_enable_data_log_force[ 891] <= 1'h0;
      write_enable_data_log_force[ 892] <= 1'h0;
      write_enable_data_log_force[ 893] <= 1'h0;
      write_enable_data_log_force[ 894] <= 1'h0;
      write_enable_data_log_force[ 895] <= 1'h0;
      write_enable_data_log_force[ 896] <= 1'h0;
      write_enable_data_log_force[ 897] <= 1'h0;
      write_enable_data_log_force[ 898] <= 1'h0;
      write_enable_data_log_force[ 899] <= 1'h0;
      write_enable_data_log_force[ 900] <= 1'h0;
      write_enable_data_log_force[ 901] <= 1'h0;
      write_enable_data_log_force[ 902] <= 1'h0;
      write_enable_data_log_force[ 903] <= 1'h0;
      write_enable_data_log_force[ 904] <= 1'h0;
      write_enable_data_log_force[ 905] <= 1'h0;
      write_enable_data_log_force[ 906] <= 1'h0;
      write_enable_data_log_force[ 907] <= 1'h0;
      write_enable_data_log_force[ 908] <= 1'h0;
      write_enable_data_log_force[ 909] <= 1'h0;
      write_enable_data_log_force[ 910] <= 1'h0;
      write_enable_data_log_force[ 911] <= 1'h0;
      write_enable_data_log_force[ 912] <= 1'h0;
      write_enable_data_log_force[ 913] <= 1'h0;
      write_enable_data_log_force[ 914] <= 1'h0;
      write_enable_data_log_force[ 915] <= 1'h0;
      write_enable_data_log_force[ 916] <= 1'h0;
      write_enable_data_log_force[ 917] <= 1'h0;
      write_enable_data_log_force[ 918] <= 1'h0;
      write_enable_data_log_force[ 919] <= 1'h0;
      write_enable_data_log_force[ 920] <= 1'h0;
      write_enable_data_log_force[ 921] <= 1'h0;
      write_enable_data_log_force[ 922] <= 1'h0;
      write_enable_data_log_force[ 923] <= 1'h0;
      write_enable_data_log_force[ 924] <= 1'h0;
      write_enable_data_log_force[ 925] <= 1'h0;
      write_enable_data_log_force[ 926] <= 1'h0;
      write_enable_data_log_force[ 927] <= 1'h0;
      write_enable_data_log_force[ 928] <= 1'h0;
      write_enable_data_log_force[ 929] <= 1'h0;
      write_enable_data_log_force[ 930] <= 1'h0;
      write_enable_data_log_force[ 931] <= 1'h0;
      write_enable_data_log_force[ 932] <= 1'h0;
      write_enable_data_log_force[ 933] <= 1'h0;
      write_enable_data_log_force[ 934] <= 1'h0;
      write_enable_data_log_force[ 935] <= 1'h0;
      write_enable_data_log_force[ 936] <= 1'h0;
      write_enable_data_log_force[ 937] <= 1'h0;
      write_enable_data_log_force[ 938] <= 1'h0;
      write_enable_data_log_force[ 939] <= 1'h0;
      write_enable_data_log_force[ 940] <= 1'h0;
      write_enable_data_log_force[ 941] <= 1'h0;
      write_enable_data_log_force[ 942] <= 1'h0;
      write_enable_data_log_force[ 943] <= 1'h0;
      write_enable_data_log_force[ 944] <= 1'h0;
      write_enable_data_log_force[ 945] <= 1'h0;
      write_enable_data_log_force[ 946] <= 1'h0;
      write_enable_data_log_force[ 947] <= 1'h0;
      write_enable_data_log_force[ 948] <= 1'h0;
      write_enable_data_log_force[ 949] <= 1'h0;
      write_enable_data_log_force[ 950] <= 1'h0;
      write_enable_data_log_force[ 951] <= 1'h0;
      write_enable_data_log_force[ 952] <= 1'h0;
      write_enable_data_log_force[ 953] <= 1'h0;
      write_enable_data_log_force[ 954] <= 1'h0;
      write_enable_data_log_force[ 955] <= 1'h0;
      write_enable_data_log_force[ 956] <= 1'h0;
      write_enable_data_log_force[ 957] <= 1'h0;
      write_enable_data_log_force[ 958] <= 1'h0;
      write_enable_data_log_force[ 959] <= 1'h0;
      write_enable_data_log_force[ 960] <= 1'h0;
      write_enable_data_log_force[ 961] <= 1'h0;
      write_enable_data_log_force[ 962] <= 1'h0;
      write_enable_data_log_force[ 963] <= 1'h0;
      write_enable_data_log_force[ 964] <= 1'h0;
      write_enable_data_log_force[ 965] <= 1'h0;
      write_enable_data_log_force[ 966] <= 1'h0;
      write_enable_data_log_force[ 967] <= 1'h0;
      write_enable_data_log_force[ 968] <= 1'h0;
      write_enable_data_log_force[ 969] <= 1'h0;
      write_enable_data_log_force[ 970] <= 1'h0;
      write_enable_data_log_force[ 971] <= 1'h0;
      write_enable_data_log_force[ 972] <= 1'h0;
      write_enable_data_log_force[ 973] <= 1'h0;
      write_enable_data_log_force[ 974] <= 1'h0;
      write_enable_data_log_force[ 975] <= 1'h0;
      write_enable_data_log_force[ 976] <= 1'h0;
      write_enable_data_log_force[ 977] <= 1'h0;
      write_enable_data_log_force[ 978] <= 1'h0;
      write_enable_data_log_force[ 979] <= 1'h0;
      write_enable_data_log_force[ 980] <= 1'h0;
      write_enable_data_log_force[ 981] <= 1'h0;
      write_enable_data_log_force[ 982] <= 1'h0;
      write_enable_data_log_force[ 983] <= 1'h0;
      write_enable_data_log_force[ 984] <= 1'h0;
      write_enable_data_log_force[ 985] <= 1'h0;
      write_enable_data_log_force[ 986] <= 1'h0;
      write_enable_data_log_force[ 987] <= 1'h0;
      write_enable_data_log_force[ 988] <= 1'h0;
      write_enable_data_log_force[ 989] <= 1'h0;
      write_enable_data_log_force[ 990] <= 1'h0;
      write_enable_data_log_force[ 991] <= 1'h0;
      write_enable_data_log_force[ 992] <= 1'h0;
      write_enable_data_log_force[ 993] <= 1'h0;
      write_enable_data_log_force[ 994] <= 1'h0;
      write_enable_data_log_force[ 995] <= 1'h0;
      write_enable_data_log_force[ 996] <= 1'h0;
      write_enable_data_log_force[ 997] <= 1'h0;
      write_enable_data_log_force[ 998] <= 1'h0;
      write_enable_data_log_force[ 999] <= 1'h0;
      write_enable_data_log_force[1000] <= 1'h0;
      write_enable_data_log_force[1001] <= 1'h0;
      write_enable_data_log_force[1002] <= 1'h0;
      write_enable_data_log_force[1003] <= 1'h0;
      write_enable_data_log_force[1004] <= 1'h0;
      write_enable_data_log_force[1005] <= 1'h0;
      write_enable_data_log_force[1006] <= 1'h0;
      write_enable_data_log_force[1007] <= 1'h0;
      write_enable_data_log_force[1008] <= 1'h0;
      write_enable_data_log_force[1009] <= 1'h0;
      write_enable_data_log_force[1010] <= 1'h0;
      write_enable_data_log_force[1011] <= 1'h0;
      write_enable_data_log_force[1012] <= 1'h0;
      write_enable_data_log_force[1013] <= 1'h0;
      write_enable_data_log_force[1014] <= 1'h0;
      write_enable_data_log_force[1015] <= 1'h0;
      write_enable_data_log_force[1016] <= 1'h0;
      write_enable_data_log_force[1017] <= 1'h0;
      write_enable_data_log_force[1018] <= 1'h0;
      write_enable_data_log_force[1019] <= 1'h0;
      write_enable_data_log_force[1020] <= 1'h0;
      write_enable_data_log_force[1021] <= 1'h0;
      write_enable_data_log_force[1022] <= 1'h0;
      write_enable_data_log_force[1023] <= 1'h0;
      write_enable_data_log_force[1024] <= 1'h0;
      write_enable_data_log_force[1025] <= 1'h0;
      write_enable_data_log_force[1026] <= 1'h0;
      write_enable_data_log_force[1027] <= 1'h0;
      write_enable_data_log_force[1028] <= 1'h0;
      write_enable_data_log_force[1029] <= 1'h0;
      write_enable_data_log_force[1030] <= 1'h0;
      write_enable_data_log_force[1031] <= 1'h0;
      write_enable_data_log_force[1032] <= 1'h0;
      write_enable_data_log_force[1033] <= 1'h0;
      write_enable_data_log_force[1034] <= 1'h0;
      write_enable_data_log_force[1035] <= 1'h0;
      write_enable_data_log_force[1036] <= 1'h0;
      write_enable_data_log_force[1037] <= 1'h0;
      write_enable_data_log_force[1038] <= 1'h0;
      write_enable_data_log_force[1039] <= 1'h0;
      write_enable_data_log_force[1040] <= 1'h0;
      write_enable_data_log_force[1041] <= 1'h0;
      write_enable_data_log_force[1042] <= 1'h0;
      write_enable_data_log_force[1043] <= 1'h0;
      write_enable_data_log_force[1044] <= 1'h0;
      write_enable_data_log_force[1045] <= 1'h0;
      write_enable_data_log_force[1046] <= 1'h0;
      write_enable_data_log_force[1047] <= 1'h0;
      write_enable_data_log_force[1048] <= 1'h0;
      write_enable_data_log_force[1049] <= 1'h0;
      write_enable_data_log_force[1050] <= 1'h0;
      write_enable_data_log_force[1051] <= 1'h0;
      write_enable_data_log_force[1052] <= 1'h0;
      write_enable_data_log_force[1053] <= 1'h0;
      write_enable_data_log_force[1054] <= 1'h0;
      write_enable_data_log_force[1055] <= 1'h0;
      write_enable_data_log_force[1056] <= 1'h0;
      write_enable_data_log_force[1057] <= 1'h0;
      write_enable_data_log_force[1058] <= 1'h0;
      write_enable_data_log_force[1059] <= 1'h0;
      write_enable_data_log_force[1060] <= 1'h0;
      write_enable_data_log_force[1061] <= 1'h0;
      write_enable_data_log_force[1062] <= 1'h0;
      write_enable_data_log_force[1063] <= 1'h0;
      write_enable_data_log_force[1064] <= 1'h0;
      write_enable_data_log_force[1065] <= 1'h0;
      write_enable_data_log_force[1066] <= 1'h0;
      write_enable_data_log_force[1067] <= 1'h0;
      write_enable_data_log_force[1068] <= 1'h0;
      write_enable_data_log_force[1069] <= 1'h0;
      write_enable_data_log_force[1070] <= 1'h0;
      write_enable_data_log_force[1071] <= 1'h0;
      write_enable_data_log_force[1072] <= 1'h0;
      write_enable_data_log_force[1073] <= 1'h0;
      write_enable_data_log_force[1074] <= 1'h0;
      write_enable_data_log_force[1075] <= 1'h0;
      write_enable_data_log_force[1076] <= 1'h0;
      write_enable_data_log_force[1077] <= 1'h0;
      write_enable_data_log_force[1078] <= 1'h0;
      write_enable_data_log_force[1079] <= 1'h0;
      write_enable_data_log_force[1080] <= 1'h0;
      write_enable_data_log_force[1081] <= 1'h0;
      write_enable_data_log_force[1082] <= 1'h0;
      write_enable_data_log_force[1083] <= 1'h0;
      write_enable_data_log_force[1084] <= 1'h0;
      write_enable_data_log_force[1085] <= 1'h0;
      write_enable_data_log_force[1086] <= 1'h0;
      write_enable_data_log_force[1087] <= 1'h0;
      write_enable_data_log_force[1088] <= 1'h0;
      write_enable_data_log_force[1089] <= 1'h0;
      write_enable_data_log_force[1090] <= 1'h0;
      write_enable_data_log_force[1091] <= 1'h0;
      write_enable_data_log_force[1092] <= 1'h0;
      write_enable_data_log_force[1093] <= 1'h0;
      write_enable_data_log_force[1094] <= 1'h0;
      write_enable_data_log_force[1095] <= 1'h0;
      write_enable_data_log_force[1096] <= 1'h0;
      write_enable_data_log_force[1097] <= 1'h0;
      write_enable_data_log_force[1098] <= 1'h0;
      write_enable_data_log_force[1099] <= 1'h0;
      write_enable_data_log_force[1100] <= 1'h0;
      write_enable_data_log_force[1101] <= 1'h0;
      write_enable_data_log_force[1102] <= 1'h0;
      write_enable_data_log_force[1103] <= 1'h0;
      write_enable_data_log_force[1104] <= 1'h0;
      write_enable_data_log_force[1105] <= 1'h0;
      write_enable_data_log_force[1106] <= 1'h0;
      write_enable_data_log_force[1107] <= 1'h0;
      write_enable_data_log_force[1108] <= 1'h0;
      write_enable_data_log_force[1109] <= 1'h0;
      write_enable_data_log_force[1110] <= 1'h0;
      write_enable_data_log_force[1111] <= 1'h0;
      write_enable_data_log_force[1112] <= 1'h0;
      write_enable_data_log_force[1113] <= 1'h0;
      write_enable_data_log_force[1114] <= 1'h0;
      write_enable_data_log_force[1115] <= 1'h0;
      write_enable_data_log_force[1116] <= 1'h0;
      write_enable_data_log_force[1117] <= 1'h0;
      write_enable_data_log_force[1118] <= 1'h0;
      write_enable_data_log_force[1119] <= 1'h0;
      write_enable_data_log_force[1120] <= 1'h0;
      write_enable_data_log_force[1121] <= 1'h0;
      write_enable_data_log_force[1122] <= 1'h0;
      write_enable_data_log_force[1123] <= 1'h0;
      write_enable_data_log_force[1124] <= 1'h0;
      write_enable_data_log_force[1125] <= 1'h0;
      write_enable_data_log_force[1126] <= 1'h0;
      write_enable_data_log_force[1127] <= 1'h0;
      write_enable_data_log_force[1128] <= 1'h0;
      write_enable_data_log_force[1129] <= 1'h0;
      write_enable_data_log_force[1130] <= 1'h0;
      write_enable_data_log_force[1131] <= 1'h0;
      write_enable_data_log_force[1132] <= 1'h0;
      write_enable_data_log_force[1133] <= 1'h0;
      write_enable_data_log_force[1134] <= 1'h0;
      write_enable_data_log_force[1135] <= 1'h0;
      write_enable_data_log_force[1136] <= 1'h0;
      write_enable_data_log_force[1137] <= 1'h0;
      write_enable_data_log_force[1138] <= 1'h0;
      write_enable_data_log_force[1139] <= 1'h0;
      write_enable_data_log_force[1140] <= 1'h0;
      write_enable_data_log_force[1141] <= 1'h0;
      write_enable_data_log_force[1142] <= 1'h0;
      write_enable_data_log_force[1143] <= 1'h0;
      write_enable_data_log_force[1144] <= 1'h0;
      write_enable_data_log_force[1145] <= 1'h0;
      write_enable_data_log_force[1146] <= 1'h0;
      write_enable_data_log_force[1147] <= 1'h0;
      write_enable_data_log_force[1148] <= 1'h0;
      write_enable_data_log_force[1149] <= 1'h0;
      write_enable_data_log_force[1150] <= 1'h0;
      write_enable_data_log_force[1151] <= 1'h0;
      write_enable_data_log_force[1152] <= 1'h0;
      write_enable_data_log_force[1153] <= 1'h0;
      write_enable_data_log_force[1154] <= 1'h0;
      write_enable_data_log_force[1155] <= 1'h0;
      write_enable_data_log_force[1156] <= 1'h0;
      write_enable_data_log_force[1157] <= 1'h0;
      write_enable_data_log_force[1158] <= 1'h0;
      write_enable_data_log_force[1159] <= 1'h0;
      write_enable_data_log_force[1160] <= 1'h0;
      write_enable_data_log_force[1161] <= 1'h0;
      write_enable_data_log_force[1162] <= 1'h0;
      write_enable_data_log_force[1163] <= 1'h0;
      write_enable_data_log_force[1164] <= 1'h0;
      write_enable_data_log_force[1165] <= 1'h0;
      write_enable_data_log_force[1166] <= 1'h0;
      write_enable_data_log_force[1167] <= 1'h0;
      write_enable_data_log_force[1168] <= 1'h0;
      write_enable_data_log_force[1169] <= 1'h0;
      write_enable_data_log_force[1170] <= 1'h0;
      write_enable_data_log_force[1171] <= 1'h0;
      write_enable_data_log_force[1172] <= 1'h0;
      write_enable_data_log_force[1173] <= 1'h0;
      write_enable_data_log_force[1174] <= 1'h0;
      write_enable_data_log_force[1175] <= 1'h0;
      write_enable_data_log_force[1176] <= 1'h0;
      write_enable_data_log_force[1177] <= 1'h0;
      write_enable_data_log_force[1178] <= 1'h0;
      write_enable_data_log_force[1179] <= 1'h0;
      write_enable_data_log_force[1180] <= 1'h0;
      write_enable_data_log_force[1181] <= 1'h0;
      write_enable_data_log_force[1182] <= 1'h0;
      write_enable_data_log_force[1183] <= 1'h0;
      write_enable_data_log_force[1184] <= 1'h0;
      write_enable_data_log_force[1185] <= 1'h0;
      write_enable_data_log_force[1186] <= 1'h0;
      write_enable_data_log_force[1187] <= 1'h0;
      write_enable_data_log_force[1188] <= 1'h0;
      write_enable_data_log_force[1189] <= 1'h0;
      write_enable_data_log_force[1190] <= 1'h0;
      write_enable_data_log_force[1191] <= 1'h0;
      write_enable_data_log_force[1192] <= 1'h0;
      write_enable_data_log_force[1193] <= 1'h0;
      write_enable_data_log_force[1194] <= 1'h0;
      write_enable_data_log_force[1195] <= 1'h0;
      write_enable_data_log_force[1196] <= 1'h0;
      write_enable_data_log_force[1197] <= 1'h0;
      write_enable_data_log_force[1198] <= 1'h0;
      write_enable_data_log_force[1199] <= 1'h0;
      write_enable_data_log_force[1200] <= 1'h0;
      write_enable_data_log_force[1201] <= 1'h0;
      write_enable_data_log_force[1202] <= 1'h0;
      write_enable_data_log_force[1203] <= 1'h0;
      write_enable_data_log_force[1204] <= 1'h0;
      write_enable_data_log_force[1205] <= 1'h0;
      write_enable_data_log_force[1206] <= 1'h0;
      write_enable_data_log_force[1207] <= 1'h0;
      write_enable_data_log_force[1208] <= 1'h0;
      write_enable_data_log_force[1209] <= 1'h0;
      write_enable_data_log_force[1210] <= 1'h0;
      write_enable_data_log_force[1211] <= 1'h0;
      write_enable_data_log_force[1212] <= 1'h0;
      write_enable_data_log_force[1213] <= 1'h0;
      write_enable_data_log_force[1214] <= 1'h0;
      write_enable_data_log_force[1215] <= 1'h0;
      write_enable_data_log_force[1216] <= 1'h0;
      write_enable_data_log_force[1217] <= 1'h0;
      write_enable_data_log_force[1218] <= 1'h0;
      write_enable_data_log_force[1219] <= 1'h0;
      write_enable_data_log_force[1220] <= 1'h0;
      write_enable_data_log_force[1221] <= 1'h0;
      write_enable_data_log_force[1222] <= 1'h0;
      write_enable_data_log_force[1223] <= 1'h0;
      write_enable_data_log_force[1224] <= 1'h0;
      write_enable_data_log_force[1225] <= 1'h0;
      write_enable_data_log_force[1226] <= 1'h0;
      write_enable_data_log_force[1227] <= 1'h0;
      write_enable_data_log_force[1228] <= 1'h0;
      write_enable_data_log_force[1229] <= 1'h0;
      write_enable_data_log_force[1230] <= 1'h0;
      write_enable_data_log_force[1231] <= 1'h0;
      write_enable_data_log_force[1232] <= 1'h0;
      write_enable_data_log_force[1233] <= 1'h0;
      write_enable_data_log_force[1234] <= 1'h0;
      write_enable_data_log_force[1235] <= 1'h0;
      write_enable_data_log_force[1236] <= 1'h0;
      write_enable_data_log_force[1237] <= 1'h0;
      write_enable_data_log_force[1238] <= 1'h0;
      write_enable_data_log_force[1239] <= 1'h0;
      write_enable_data_log_force[1240] <= 1'h0;
      write_enable_data_log_force[1241] <= 1'h0;
      write_enable_data_log_force[1242] <= 1'h0;
      write_enable_data_log_force[1243] <= 1'h0;
      write_enable_data_log_force[1244] <= 1'h0;
      write_enable_data_log_force[1245] <= 1'h0;
      write_enable_data_log_force[1246] <= 1'h0;
      write_enable_data_log_force[1247] <= 1'h0;
      write_enable_data_log_force[1248] <= 1'h0;
      write_enable_data_log_force[1249] <= 1'h0;
      write_enable_data_log_force[1250] <= 1'h0;
      write_enable_data_log_force[1251] <= 1'h0;
      write_enable_data_log_force[1252] <= 1'h0;
      write_enable_data_log_force[1253] <= 1'h0;
      write_enable_data_log_force[1254] <= 1'h0;
      write_enable_data_log_force[1255] <= 1'h0;
      write_enable_data_log_force[1256] <= 1'h0;
      write_enable_data_log_force[1257] <= 1'h0;
      write_enable_data_log_force[1258] <= 1'h0;
      write_enable_data_log_force[1259] <= 1'h0;
      write_enable_data_log_force[1260] <= 1'h0;
      write_enable_data_log_force[1261] <= 1'h0;
      write_enable_data_log_force[1262] <= 1'h0;
      write_enable_data_log_force[1263] <= 1'h0;
      write_enable_data_log_force[1264] <= 1'h0;
      write_enable_data_log_force[1265] <= 1'h0;
      write_enable_data_log_force[1266] <= 1'h0;
      write_enable_data_log_force[1267] <= 1'h0;
      write_enable_data_log_force[1268] <= 1'h0;
      write_enable_data_log_force[1269] <= 1'h0;
      write_enable_data_log_force[1270] <= 1'h0;
      write_enable_data_log_force[1271] <= 1'h0;
      write_enable_data_log_force[1272] <= 1'h0;
      write_enable_data_log_force[1273] <= 1'h0;
      write_enable_data_log_force[1274] <= 1'h0;
      write_enable_data_log_force[1275] <= 1'h0;
      write_enable_data_log_force[1276] <= 1'h0;
      write_enable_data_log_force[1277] <= 1'h0;
      write_enable_data_log_force[1278] <= 1'h0;
      write_enable_data_log_force[1279] <= 1'h0;
      write_enable_data_log_force[1280] <= 1'h0;
      write_enable_data_log_force[1281] <= 1'h0;
      write_enable_data_log_force[1282] <= 1'h0;
      write_enable_data_log_force[1283] <= 1'h0;
      write_enable_data_log_force[1284] <= 1'h0;
      write_enable_data_log_force[1285] <= 1'h0;
      write_enable_data_log_force[1286] <= 1'h0;
      write_enable_data_log_force[1287] <= 1'h0;
      write_enable_data_log_force[1288] <= 1'h0;
      write_enable_data_log_force[1289] <= 1'h0;
      write_enable_data_log_force[1290] <= 1'h0;
      write_enable_data_log_force[1291] <= 1'h0;
      write_enable_data_log_force[1292] <= 1'h0;
      write_enable_data_log_force[1293] <= 1'h0;
      write_enable_data_log_force[1294] <= 1'h0;
      write_enable_data_log_force[1295] <= 1'h0;
      write_enable_data_log_force[1296] <= 1'h0;
      write_enable_data_log_force[1297] <= 1'h0;
      write_enable_data_log_force[1298] <= 1'h0;
      write_enable_data_log_force[1299] <= 1'h0;
      write_enable_data_log_force[1300] <= 1'h0;
      write_enable_data_log_force[1301] <= 1'h0;
      write_enable_data_log_force[1302] <= 1'h0;
      write_enable_data_log_force[1303] <= 1'h0;
      write_enable_data_log_force[1304] <= 1'h0;
      write_enable_data_log_force[1305] <= 1'h0;
      write_enable_data_log_force[1306] <= 1'h0;
      write_enable_data_log_force[1307] <= 1'h0;
      write_enable_data_log_force[1308] <= 1'h0;
      write_enable_data_log_force[1309] <= 1'h0;
      write_enable_data_log_force[1310] <= 1'h0;
      write_enable_data_log_force[1311] <= 1'h0;
      write_enable_data_log_force[1312] <= 1'h0;
      write_enable_data_log_force[1313] <= 1'h0;
      write_enable_data_log_force[1314] <= 1'h0;
      write_enable_data_log_force[1315] <= 1'h0;
      write_enable_data_log_force[1316] <= 1'h0;
      write_enable_data_log_force[1317] <= 1'h0;
      write_enable_data_log_force[1318] <= 1'h0;
      write_enable_data_log_force[1319] <= 1'h0;
      write_enable_data_log_force[1320] <= 1'h0;
      write_enable_data_log_force[1321] <= 1'h0;
      write_enable_data_log_force[1322] <= 1'h0;
      write_enable_data_log_force[1323] <= 1'h0;
      write_enable_data_log_force[1324] <= 1'h0;
      write_enable_data_log_force[1325] <= 1'h0;
      write_enable_data_log_force[1326] <= 1'h0;
      write_enable_data_log_force[1327] <= 1'h0;
      write_enable_data_log_force[1328] <= 1'h0;
      write_enable_data_log_force[1329] <= 1'h0;
      write_enable_data_log_force[1330] <= 1'h0;
      write_enable_data_log_force[1331] <= 1'h0;
      write_enable_data_log_force[1332] <= 1'h0;
      write_enable_data_log_force[1333] <= 1'h0;
      write_enable_data_log_force[1334] <= 1'h0;
      write_enable_data_log_force[1335] <= 1'h0;
      write_enable_data_log_force[1336] <= 1'h0;
      write_enable_data_log_force[1337] <= 1'h0;
      write_enable_data_log_force[1338] <= 1'h0;
      write_enable_data_log_force[1339] <= 1'h0;
      write_enable_data_log_force[1340] <= 1'h0;
      write_enable_data_log_force[1341] <= 1'h0;
      write_enable_data_log_force[1342] <= 1'h0;
      write_enable_data_log_force[1343] <= 1'h0;
      write_enable_data_log_force[1344] <= 1'h0;
      write_enable_data_log_force[1345] <= 1'h0;
      write_enable_data_log_force[1346] <= 1'h0;
      write_enable_data_log_force[1347] <= 1'h0;
      write_enable_data_log_force[1348] <= 1'h0;
      write_enable_data_log_force[1349] <= 1'h0;
      write_enable_data_log_force[1350] <= 1'h0;
      write_enable_data_log_force[1351] <= 1'h0;
      write_enable_data_log_force[1352] <= 1'h0;
      write_enable_data_log_force[1353] <= 1'h0;
      write_enable_data_log_force[1354] <= 1'h0;
      write_enable_data_log_force[1355] <= 1'h0;
      write_enable_data_log_force[1356] <= 1'h0;
      write_enable_data_log_force[1357] <= 1'h0;
      write_enable_data_log_force[1358] <= 1'h0;
      write_enable_data_log_force[1359] <= 1'h0;
      write_enable_data_log_force[1360] <= 1'h0;
      write_enable_data_log_force[1361] <= 1'h0;
      write_enable_data_log_force[1362] <= 1'h0;
      write_enable_data_log_force[1363] <= 1'h0;
      write_enable_data_log_force[1364] <= 1'h0;
      write_enable_data_log_force[1365] <= 1'h0;
      write_enable_data_log_force[1366] <= 1'h0;
      write_enable_data_log_force[1367] <= 1'h0;
      write_enable_data_log_force[1368] <= 1'h0;
      write_enable_data_log_force[1369] <= 1'h0;
      write_enable_data_log_force[1370] <= 1'h0;
      write_enable_data_log_force[1371] <= 1'h0;
      write_enable_data_log_force[1372] <= 1'h0;
      write_enable_data_log_force[1373] <= 1'h0;
      write_enable_data_log_force[1374] <= 1'h0;
      write_enable_data_log_force[1375] <= 1'h0;
      write_enable_data_log_force[1376] <= 1'h0;
      write_enable_data_log_force[1377] <= 1'h0;
      write_enable_data_log_force[1378] <= 1'h0;
      write_enable_data_log_force[1379] <= 1'h0;
      write_enable_data_log_force[1380] <= 1'h0;
      write_enable_data_log_force[1381] <= 1'h0;
      write_enable_data_log_force[1382] <= 1'h0;
      write_enable_data_log_force[1383] <= 1'h0;
      write_enable_data_log_force[1384] <= 1'h0;
      write_enable_data_log_force[1385] <= 1'h0;
      write_enable_data_log_force[1386] <= 1'h0;
      write_enable_data_log_force[1387] <= 1'h0;
      write_enable_data_log_force[1388] <= 1'h0;
      write_enable_data_log_force[1389] <= 1'h0;
      write_enable_data_log_force[1390] <= 1'h0;
      write_enable_data_log_force[1391] <= 1'h0;
      write_enable_data_log_force[1392] <= 1'h0;
      write_enable_data_log_force[1393] <= 1'h0;
      write_enable_data_log_force[1394] <= 1'h0;
      write_enable_data_log_force[1395] <= 1'h0;
      write_enable_data_log_force[1396] <= 1'h0;
      write_enable_data_log_force[1397] <= 1'h0;
      write_enable_data_log_force[1398] <= 1'h0;
      write_enable_data_log_force[1399] <= 1'h0;
      write_enable_data_log_force[1400] <= 1'h0;
      write_enable_data_log_force[1401] <= 1'h0;
      write_enable_data_log_force[1402] <= 1'h0;
      write_enable_data_log_force[1403] <= 1'h0;
      write_enable_data_log_force[1404] <= 1'h0;
      write_enable_data_log_force[1405] <= 1'h0;
      write_enable_data_log_force[1406] <= 1'h0;
      write_enable_data_log_force[1407] <= 1'h0;
      write_enable_data_log_force[1408] <= 1'h0;
      write_enable_data_log_force[1409] <= 1'h0;
      write_enable_data_log_force[1410] <= 1'h0;
      write_enable_data_log_force[1411] <= 1'h0;
      write_enable_data_log_force[1412] <= 1'h0;
      write_enable_data_log_force[1413] <= 1'h0;
      write_enable_data_log_force[1414] <= 1'h0;
      write_enable_data_log_force[1415] <= 1'h0;
      write_enable_data_log_force[1416] <= 1'h0;
      write_enable_data_log_force[1417] <= 1'h0;
      write_enable_data_log_force[1418] <= 1'h0;
      write_enable_data_log_force[1419] <= 1'h0;
      write_enable_data_log_force[1420] <= 1'h0;
      write_enable_data_log_force[1421] <= 1'h0;
      write_enable_data_log_force[1422] <= 1'h0;
      write_enable_data_log_force[1423] <= 1'h0;
      write_enable_data_log_force[1424] <= 1'h0;
      write_enable_data_log_force[1425] <= 1'h0;
      write_enable_data_log_force[1426] <= 1'h0;
      write_enable_data_log_force[1427] <= 1'h0;
      write_enable_data_log_force[1428] <= 1'h0;
      write_enable_data_log_force[1429] <= 1'h0;
      write_enable_data_log_force[1430] <= 1'h0;
      write_enable_data_log_force[1431] <= 1'h0;
      write_enable_data_log_force[1432] <= 1'h0;
      write_enable_data_log_force[1433] <= 1'h0;
      write_enable_data_log_force[1434] <= 1'h0;
      write_enable_data_log_force[1435] <= 1'h0;
      write_enable_data_log_force[1436] <= 1'h0;
      write_enable_data_log_force[1437] <= 1'h0;
      write_enable_data_log_force[1438] <= 1'h0;
      write_enable_data_log_force[1439] <= 1'h0;
      write_enable_data_log_force[1440] <= 1'h0;
      write_enable_data_log_force[1441] <= 1'h0;
      write_enable_data_log_force[1442] <= 1'h0;
      write_enable_data_log_force[1443] <= 1'h0;
      write_enable_data_log_force[1444] <= 1'h0;
      write_enable_data_log_force[1445] <= 1'h0;
      write_enable_data_log_force[1446] <= 1'h0;
      write_enable_data_log_force[1447] <= 1'h0;
      write_enable_data_log_force[1448] <= 1'h0;
      write_enable_data_log_force[1449] <= 1'h0;
      write_enable_data_log_force[1450] <= 1'h0;
      write_enable_data_log_force[1451] <= 1'h0;
      write_enable_data_log_force[1452] <= 1'h0;
      write_enable_data_log_force[1453] <= 1'h0;
      write_enable_data_log_force[1454] <= 1'h0;
      write_enable_data_log_force[1455] <= 1'h0;
      write_enable_data_log_force[1456] <= 1'h0;
      write_enable_data_log_force[1457] <= 1'h0;
      write_enable_data_log_force[1458] <= 1'h0;
      write_enable_data_log_force[1459] <= 1'h0;
      write_enable_data_log_force[1460] <= 1'h0;
      write_enable_data_log_force[1461] <= 1'h0;
      write_enable_data_log_force[1462] <= 1'h0;
      write_enable_data_log_force[1463] <= 1'h0;
      write_enable_data_log_force[1464] <= 1'h0;
      write_enable_data_log_force[1465] <= 1'h0;
      write_enable_data_log_force[1466] <= 1'h0;
      write_enable_data_log_force[1467] <= 1'h0;
      write_enable_data_log_force[1468] <= 1'h0;
      write_enable_data_log_force[1469] <= 1'h0;
      write_enable_data_log_force[1470] <= 1'h0;
      write_enable_data_log_force[1471] <= 1'h0;
      write_enable_data_log_force[1472] <= 1'h0;
      write_enable_data_log_force[1473] <= 1'h0;
      write_enable_data_log_force[1474] <= 1'h0;
      write_enable_data_log_force[1475] <= 1'h0;
      write_enable_data_log_force[1476] <= 1'h0;
      write_enable_data_log_force[1477] <= 1'h0;
      write_enable_data_log_force[1478] <= 1'h0;
      write_enable_data_log_force[1479] <= 1'h0;
      write_enable_data_log_force[1480] <= 1'h0;
      write_enable_data_log_force[1481] <= 1'h0;
      write_enable_data_log_force[1482] <= 1'h0;
      write_enable_data_log_force[1483] <= 1'h0;
      write_enable_data_log_force[1484] <= 1'h0;
      write_enable_data_log_force[1485] <= 1'h0;
      write_enable_data_log_force[1486] <= 1'h0;
      write_enable_data_log_force[1487] <= 1'h0;
      write_enable_data_log_force[1488] <= 1'h0;
      write_enable_data_log_force[1489] <= 1'h0;
      write_enable_data_log_force[1490] <= 1'h0;
      write_enable_data_log_force[1491] <= 1'h0;
      write_enable_data_log_force[1492] <= 1'h0;
      write_enable_data_log_force[1493] <= 1'h0;
      write_enable_data_log_force[1494] <= 1'h0;
      write_enable_data_log_force[1495] <= 1'h0;
      write_enable_data_log_force[1496] <= 1'h0;
      write_enable_data_log_force[1497] <= 1'h0;
      write_enable_data_log_force[1498] <= 1'h0;
      write_enable_data_log_force[1499] <= 1'h0;
      write_enable_data_log_force[1500] <= 1'h0;
      write_enable_data_log_force[1501] <= 1'h0;
      write_enable_data_log_force[1502] <= 1'h0;
      write_enable_data_log_force[1503] <= 1'h0;
      write_enable_data_log_force[1504] <= 1'h0;
      write_enable_data_log_force[1505] <= 1'h0;
      write_enable_data_log_force[1506] <= 1'h0;
      write_enable_data_log_force[1507] <= 1'h0;
      write_enable_data_log_force[1508] <= 1'h0;
      write_enable_data_log_force[1509] <= 1'h0;
      write_enable_data_log_force[1510] <= 1'h0;
      write_enable_data_log_force[1511] <= 1'h0;
      write_enable_data_log_force[1512] <= 1'h0;
      write_enable_data_log_force[1513] <= 1'h0;
      write_enable_data_log_force[1514] <= 1'h0;
      write_enable_data_log_force[1515] <= 1'h0;
      write_enable_data_log_force[1516] <= 1'h0;
      write_enable_data_log_force[1517] <= 1'h0;
      write_enable_data_log_force[1518] <= 1'h0;
      write_enable_data_log_force[1519] <= 1'h0;
      write_enable_data_log_force[1520] <= 1'h0;
      write_enable_data_log_force[1521] <= 1'h0;
      write_enable_data_log_force[1522] <= 1'h0;
      write_enable_data_log_force[1523] <= 1'h0;
      write_enable_data_log_force[1524] <= 1'h0;
      write_enable_data_log_force[1525] <= 1'h0;
      write_enable_data_log_force[1526] <= 1'h0;
      write_enable_data_log_force[1527] <= 1'h0;
      write_enable_data_log_force[1528] <= 1'h0;
      write_enable_data_log_force[1529] <= 1'h0;
      write_enable_data_log_force[1530] <= 1'h0;
      write_enable_data_log_force[1531] <= 1'h0;
      write_enable_data_log_force[1532] <= 1'h0;
      write_enable_data_log_force[1533] <= 1'h0;
      write_enable_data_log_force[1534] <= 1'h0;
      write_enable_data_log_force[1535] <= 1'h0;
      write_enable_data_log_force[1536] <= 1'h0;
      write_enable_data_log_force[1537] <= 1'h0;
      write_enable_data_log_force[1538] <= 1'h0;
      write_enable_data_log_force[1539] <= 1'h0;
      write_enable_data_log_force[1540] <= 1'h0;
      write_enable_data_log_force[1541] <= 1'h0;
      write_enable_data_log_force[1542] <= 1'h0;
      write_enable_data_log_force[1543] <= 1'h0;
      write_enable_data_log_force[1544] <= 1'h0;
      write_enable_data_log_force[1545] <= 1'h0;
      write_enable_data_log_force[1546] <= 1'h0;
      write_enable_data_log_force[1547] <= 1'h0;
      write_enable_data_log_force[1548] <= 1'h0;
      write_enable_data_log_force[1549] <= 1'h0;
      write_enable_data_log_force[1550] <= 1'h0;
      write_enable_data_log_force[1551] <= 1'h0;
      write_enable_data_log_force[1552] <= 1'h0;
      write_enable_data_log_force[1553] <= 1'h0;
      write_enable_data_log_force[1554] <= 1'h0;
      write_enable_data_log_force[1555] <= 1'h0;
      write_enable_data_log_force[1556] <= 1'h0;
      write_enable_data_log_force[1557] <= 1'h0;
      write_enable_data_log_force[1558] <= 1'h0;
      write_enable_data_log_force[1559] <= 1'h0;
      write_enable_data_log_force[1560] <= 1'h0;
      write_enable_data_log_force[1561] <= 1'h0;
      write_enable_data_log_force[1562] <= 1'h0;
      write_enable_data_log_force[1563] <= 1'h0;
      write_enable_data_log_force[1564] <= 1'h0;
      write_enable_data_log_force[1565] <= 1'h0;
      write_enable_data_log_force[1566] <= 1'h0;
      write_enable_data_log_force[1567] <= 1'h0;
      write_enable_data_log_force[1568] <= 1'h0;
      write_enable_data_log_force[1569] <= 1'h0;
      write_enable_data_log_force[1570] <= 1'h0;
      write_enable_data_log_force[1571] <= 1'h0;
      write_enable_data_log_force[1572] <= 1'h0;
      write_enable_data_log_force[1573] <= 1'h0;
      write_enable_data_log_force[1574] <= 1'h0;
      write_enable_data_log_force[1575] <= 1'h0;
      write_enable_data_log_force[1576] <= 1'h0;
      write_enable_data_log_force[1577] <= 1'h0;
      write_enable_data_log_force[1578] <= 1'h0;
      write_enable_data_log_force[1579] <= 1'h0;
      write_enable_data_log_force[1580] <= 1'h0;
      write_enable_data_log_force[1581] <= 1'h0;
      write_enable_data_log_force[1582] <= 1'h0;
      write_enable_data_log_force[1583] <= 1'h0;
      write_enable_data_log_force[1584] <= 1'h0;
      write_enable_data_log_force[1585] <= 1'h0;
      write_enable_data_log_force[1586] <= 1'h0;
      write_enable_data_log_force[1587] <= 1'h0;
      write_enable_data_log_force[1588] <= 1'h0;
      write_enable_data_log_force[1589] <= 1'h0;
      write_enable_data_log_force[1590] <= 1'h0;
      write_enable_data_log_force[1591] <= 1'h0;
      write_enable_data_log_force[1592] <= 1'h0;
      write_enable_data_log_force[1593] <= 1'h0;
      write_enable_data_log_force[1594] <= 1'h0;
      write_enable_data_log_force[1595] <= 1'h0;
      write_enable_data_log_force[1596] <= 1'h0;
      write_enable_data_log_force[1597] <= 1'h0;
      write_enable_data_log_force[1598] <= 1'h0;
      write_enable_data_log_force[1599] <= 1'h0;
      write_enable_data_log_force[1600] <= 1'h0;
      write_enable_data_log_force[1601] <= 1'h0;
      write_enable_data_log_force[1602] <= 1'h0;
      write_enable_data_log_force[1603] <= 1'h0;
      write_enable_data_log_force[1604] <= 1'h0;
      write_enable_data_log_force[1605] <= 1'h0;
      write_enable_data_log_force[1606] <= 1'h0;
      write_enable_data_log_force[1607] <= 1'h0;
      write_enable_data_log_force[1608] <= 1'h0;
      write_enable_data_log_force[1609] <= 1'h0;
      write_enable_data_log_force[1610] <= 1'h0;
      write_enable_data_log_force[1611] <= 1'h0;
      write_enable_data_log_force[1612] <= 1'h0;
      write_enable_data_log_force[1613] <= 1'h0;
      write_enable_data_log_force[1614] <= 1'h0;
      write_enable_data_log_force[1615] <= 1'h0;
      write_enable_data_log_force[1616] <= 1'h0;
      write_enable_data_log_force[1617] <= 1'h0;
      write_enable_data_log_force[1618] <= 1'h0;
      write_enable_data_log_force[1619] <= 1'h0;
      write_enable_data_log_force[1620] <= 1'h0;
      write_enable_data_log_force[1621] <= 1'h0;
      write_enable_data_log_force[1622] <= 1'h0;
      write_enable_data_log_force[1623] <= 1'h0;
      write_enable_data_log_force[1624] <= 1'h0;
      write_enable_data_log_force[1625] <= 1'h0;
      write_enable_data_log_force[1626] <= 1'h0;
      write_enable_data_log_force[1627] <= 1'h0;
      write_enable_data_log_force[1628] <= 1'h0;
      write_enable_data_log_force[1629] <= 1'h0;
      write_enable_data_log_force[1630] <= 1'h0;
      write_enable_data_log_force[1631] <= 1'h0;
      write_enable_data_log_force[1632] <= 1'h0;
      write_enable_data_log_force[1633] <= 1'h0;
      write_enable_data_log_force[1634] <= 1'h0;
      write_enable_data_log_force[1635] <= 1'h0;
      write_enable_data_log_force[1636] <= 1'h0;
      write_enable_data_log_force[1637] <= 1'h0;
      write_enable_data_log_force[1638] <= 1'h0;
      write_enable_data_log_force[1639] <= 1'h0;
      write_enable_data_log_force[1640] <= 1'h0;
      write_enable_data_log_force[1641] <= 1'h0;
      write_enable_data_log_force[1642] <= 1'h0;
      write_enable_data_log_force[1643] <= 1'h0;
      write_enable_data_log_force[1644] <= 1'h0;
      write_enable_data_log_force[1645] <= 1'h0;
      write_enable_data_log_force[1646] <= 1'h0;
      write_enable_data_log_force[1647] <= 1'h0;
      write_enable_data_log_force[1648] <= 1'h0;
      write_enable_data_log_force[1649] <= 1'h0;
      write_enable_data_log_force[1650] <= 1'h0;
      write_enable_data_log_force[1651] <= 1'h0;
      write_enable_data_log_force[1652] <= 1'h0;
      write_enable_data_log_force[1653] <= 1'h0;
      write_enable_data_log_force[1654] <= 1'h0;
      write_enable_data_log_force[1655] <= 1'h0;
      write_enable_data_log_force[1656] <= 1'h0;
      write_enable_data_log_force[1657] <= 1'h0;
      write_enable_data_log_force[1658] <= 1'h0;
      write_enable_data_log_force[1659] <= 1'h0;
      write_enable_data_log_force[1660] <= 1'h0;
      write_enable_data_log_force[1661] <= 1'h0;
      write_enable_data_log_force[1662] <= 1'h0;
      write_enable_data_log_force[1663] <= 1'h0;
      write_enable_data_log_force[1664] <= 1'h0;
      write_enable_data_log_force[1665] <= 1'h0;
      write_enable_data_log_force[1666] <= 1'h0;
      write_enable_data_log_force[1667] <= 1'h0;
      write_enable_data_log_force[1668] <= 1'h0;
      write_enable_data_log_force[1669] <= 1'h0;
      write_enable_data_log_force[1670] <= 1'h0;
      write_enable_data_log_force[1671] <= 1'h0;
      write_enable_data_log_force[1672] <= 1'h0;
      write_enable_data_log_force[1673] <= 1'h0;
      write_enable_data_log_force[1674] <= 1'h0;
      write_enable_data_log_force[1675] <= 1'h0;
      write_enable_data_log_force[1676] <= 1'h0;
      write_enable_data_log_force[1677] <= 1'h0;
      write_enable_data_log_force[1678] <= 1'h0;
      write_enable_data_log_force[1679] <= 1'h0;
      write_enable_data_log_force[1680] <= 1'h0;
      write_enable_data_log_force[1681] <= 1'h0;
      write_enable_data_log_force[1682] <= 1'h0;
      write_enable_data_log_force[1683] <= 1'h0;
      write_enable_data_log_force[1684] <= 1'h0;
      write_enable_data_log_force[1685] <= 1'h0;
      write_enable_data_log_force[1686] <= 1'h0;
      write_enable_data_log_force[1687] <= 1'h0;
      write_enable_data_log_force[1688] <= 1'h0;
      write_enable_data_log_force[1689] <= 1'h0;
      write_enable_data_log_force[1690] <= 1'h0;
      write_enable_data_log_force[1691] <= 1'h0;
      write_enable_data_log_force[1692] <= 1'h0;
      write_enable_data_log_force[1693] <= 1'h0;
      write_enable_data_log_force[1694] <= 1'h0;
      write_enable_data_log_force[1695] <= 1'h0;
      write_enable_data_log_force[1696] <= 1'h0;
      write_enable_data_log_force[1697] <= 1'h0;
      write_enable_data_log_force[1698] <= 1'h0;
      write_enable_data_log_force[1699] <= 1'h0;
      write_enable_data_log_force[1700] <= 1'h0;
      write_enable_data_log_force[1701] <= 1'h0;
      write_enable_data_log_force[1702] <= 1'h0;
      write_enable_data_log_force[1703] <= 1'h0;
      write_enable_data_log_force[1704] <= 1'h0;
      write_enable_data_log_force[1705] <= 1'h0;
      write_enable_data_log_force[1706] <= 1'h0;
      write_enable_data_log_force[1707] <= 1'h0;
      write_enable_data_log_force[1708] <= 1'h0;
      write_enable_data_log_force[1709] <= 1'h0;
      write_enable_data_log_force[1710] <= 1'h0;
      write_enable_data_log_force[1711] <= 1'h0;
      write_enable_data_log_force[1712] <= 1'h0;
      write_enable_data_log_force[1713] <= 1'h0;
      write_enable_data_log_force[1714] <= 1'h0;
      write_enable_data_log_force[1715] <= 1'h0;
      write_enable_data_log_force[1716] <= 1'h0;
      write_enable_data_log_force[1717] <= 1'h0;
      write_enable_data_log_force[1718] <= 1'h0;
      write_enable_data_log_force[1719] <= 1'h0;
      write_enable_data_log_force[1720] <= 1'h0;
      write_enable_data_log_force[1721] <= 1'h0;
      write_enable_data_log_force[1722] <= 1'h0;
      write_enable_data_log_force[1723] <= 1'h0;
      write_enable_data_log_force[1724] <= 1'h0;
      write_enable_data_log_force[1725] <= 1'h0;
      write_enable_data_log_force[1726] <= 1'h0;
      write_enable_data_log_force[1727] <= 1'h0;
      write_enable_data_log_force[1728] <= 1'h0;
      write_enable_data_log_force[1729] <= 1'h0;
      write_enable_data_log_force[1730] <= 1'h0;
      write_enable_data_log_force[1731] <= 1'h0;
      write_enable_data_log_force[1732] <= 1'h0;
      write_enable_data_log_force[1733] <= 1'h0;
      write_enable_data_log_force[1734] <= 1'h0;
      write_enable_data_log_force[1735] <= 1'h0;
      write_enable_data_log_force[1736] <= 1'h0;
      write_enable_data_log_force[1737] <= 1'h0;
      write_enable_data_log_force[1738] <= 1'h0;
      write_enable_data_log_force[1739] <= 1'h0;
      write_enable_data_log_force[1740] <= 1'h0;
      write_enable_data_log_force[1741] <= 1'h0;
      write_enable_data_log_force[1742] <= 1'h0;
      write_enable_data_log_force[1743] <= 1'h0;
      write_enable_data_log_force[1744] <= 1'h0;
      write_enable_data_log_force[1745] <= 1'h0;
      write_enable_data_log_force[1746] <= 1'h0;
      write_enable_data_log_force[1747] <= 1'h0;
      write_enable_data_log_force[1748] <= 1'h0;
      write_enable_data_log_force[1749] <= 1'h0;
      write_enable_data_log_force[1750] <= 1'h0;
      write_enable_data_log_force[1751] <= 1'h0;
      write_enable_data_log_force[1752] <= 1'h0;
      write_enable_data_log_force[1753] <= 1'h0;
      write_enable_data_log_force[1754] <= 1'h0;
      write_enable_data_log_force[1755] <= 1'h0;
      write_enable_data_log_force[1756] <= 1'h0;
      write_enable_data_log_force[1757] <= 1'h0;
      write_enable_data_log_force[1758] <= 1'h0;
      write_enable_data_log_force[1759] <= 1'h0;
      write_enable_data_log_force[1760] <= 1'h0;
      write_enable_data_log_force[1761] <= 1'h0;
      write_enable_data_log_force[1762] <= 1'h0;
      write_enable_data_log_force[1763] <= 1'h0;
      write_enable_data_log_force[1764] <= 1'h0;
      write_enable_data_log_force[1765] <= 1'h0;
      write_enable_data_log_force[1766] <= 1'h0;
      write_enable_data_log_force[1767] <= 1'h0;
      write_enable_data_log_force[1768] <= 1'h0;
      write_enable_data_log_force[1769] <= 1'h0;
      write_enable_data_log_force[1770] <= 1'h0;
      write_enable_data_log_force[1771] <= 1'h0;
      write_enable_data_log_force[1772] <= 1'h0;
      write_enable_data_log_force[1773] <= 1'h0;
      write_enable_data_log_force[1774] <= 1'h0;
      write_enable_data_log_force[1775] <= 1'h0;
      write_enable_data_log_force[1776] <= 1'h0;
      write_enable_data_log_force[1777] <= 1'h0;
      write_enable_data_log_force[1778] <= 1'h0;
      write_enable_data_log_force[1779] <= 1'h0;
      write_enable_data_log_force[1780] <= 1'h0;
      write_enable_data_log_force[1781] <= 1'h0;
      write_enable_data_log_force[1782] <= 1'h0;
      write_enable_data_log_force[1783] <= 1'h0;
      write_enable_data_log_force[1784] <= 1'h0;
      write_enable_data_log_force[1785] <= 1'h0;
      write_enable_data_log_force[1786] <= 1'h0;
      write_enable_data_log_force[1787] <= 1'h0;
      write_enable_data_log_force[1788] <= 1'h0;
      write_enable_data_log_force[1789] <= 1'h0;
      write_enable_data_log_force[1790] <= 1'h0;
      write_enable_data_log_force[1791] <= 1'h0;
      write_enable_data_log_force[1792] <= 1'h0;
      write_enable_data_log_force[1793] <= 1'h0;
      write_enable_data_log_force[1794] <= 1'h0;
      write_enable_data_log_force[1795] <= 1'h0;
      write_enable_data_log_force[1796] <= 1'h0;
      write_enable_data_log_force[1797] <= 1'h0;
      write_enable_data_log_force[1798] <= 1'h0;
      write_enable_data_log_force[1799] <= 1'h0;
      write_enable_data_log_force[1800] <= 1'h0;
      write_enable_data_log_force[1801] <= 1'h0;
      write_enable_data_log_force[1802] <= 1'h0;
      write_enable_data_log_force[1803] <= 1'h0;
      write_enable_data_log_force[1804] <= 1'h0;
      write_enable_data_log_force[1805] <= 1'h0;
      write_enable_data_log_force[1806] <= 1'h0;
      write_enable_data_log_force[1807] <= 1'h0;
      write_enable_data_log_force[1808] <= 1'h0;
      write_enable_data_log_force[1809] <= 1'h0;
      write_enable_data_log_force[1810] <= 1'h0;
      write_enable_data_log_force[1811] <= 1'h0;
      write_enable_data_log_force[1812] <= 1'h0;
      write_enable_data_log_force[1813] <= 1'h0;
      write_enable_data_log_force[1814] <= 1'h0;
      write_enable_data_log_force[1815] <= 1'h0;
      write_enable_data_log_force[1816] <= 1'h0;
      write_enable_data_log_force[1817] <= 1'h0;
      write_enable_data_log_force[1818] <= 1'h0;
      write_enable_data_log_force[1819] <= 1'h0;
      write_enable_data_log_force[1820] <= 1'h0;
      write_enable_data_log_force[1821] <= 1'h0;
      write_enable_data_log_force[1822] <= 1'h0;
      write_enable_data_log_force[1823] <= 1'h0;
      write_enable_data_log_force[1824] <= 1'h0;
      write_enable_data_log_force[1825] <= 1'h0;
      write_enable_data_log_force[1826] <= 1'h0;
      write_enable_data_log_force[1827] <= 1'h0;
      write_enable_data_log_force[1828] <= 1'h0;
      write_enable_data_log_force[1829] <= 1'h0;
      write_enable_data_log_force[1830] <= 1'h0;
      write_enable_data_log_force[1831] <= 1'h0;
      write_enable_data_log_force[1832] <= 1'h0;
      write_enable_data_log_force[1833] <= 1'h0;
      write_enable_data_log_force[1834] <= 1'h0;
      write_enable_data_log_force[1835] <= 1'h0;
      write_enable_data_log_force[1836] <= 1'h0;
      write_enable_data_log_force[1837] <= 1'h0;
      write_enable_data_log_force[1838] <= 1'h0;
      write_enable_data_log_force[1839] <= 1'h0;
      write_enable_data_log_force[1840] <= 1'h0;
      write_enable_data_log_force[1841] <= 1'h0;
      write_enable_data_log_force[1842] <= 1'h0;
      write_enable_data_log_force[1843] <= 1'h0;
      write_enable_data_log_force[1844] <= 1'h0;
      write_enable_data_log_force[1845] <= 1'h0;
      write_enable_data_log_force[1846] <= 1'h0;
      write_enable_data_log_force[1847] <= 1'h0;
      write_enable_data_log_force[1848] <= 1'h0;
      write_enable_data_log_force[1849] <= 1'h0;
      write_enable_data_log_force[1850] <= 1'h0;
      write_enable_data_log_force[1851] <= 1'h0;
      write_enable_data_log_force[1852] <= 1'h0;
      write_enable_data_log_force[1853] <= 1'h0;
      write_enable_data_log_force[1854] <= 1'h0;
      write_enable_data_log_force[1855] <= 1'h0;
      write_enable_data_log_force[1856] <= 1'h0;
      write_enable_data_log_force[1857] <= 1'h0;
      write_enable_data_log_force[1858] <= 1'h0;
      write_enable_data_log_force[1859] <= 1'h0;
      write_enable_data_log_force[1860] <= 1'h0;
      write_enable_data_log_force[1861] <= 1'h0;
      write_enable_data_log_force[1862] <= 1'h0;
      write_enable_data_log_force[1863] <= 1'h0;
      write_enable_data_log_force[1864] <= 1'h0;
      write_enable_data_log_force[1865] <= 1'h0;
      write_enable_data_log_force[1866] <= 1'h0;
      write_enable_data_log_force[1867] <= 1'h0;
      write_enable_data_log_force[1868] <= 1'h0;
      write_enable_data_log_force[1869] <= 1'h0;
      write_enable_data_log_force[1870] <= 1'h0;
      write_enable_data_log_force[1871] <= 1'h0;
      write_enable_data_log_force[1872] <= 1'h0;
      write_enable_data_log_force[1873] <= 1'h0;
      write_enable_data_log_force[1874] <= 1'h0;
      write_enable_data_log_force[1875] <= 1'h0;
      write_enable_data_log_force[1876] <= 1'h0;
      write_enable_data_log_force[1877] <= 1'h0;
      write_enable_data_log_force[1878] <= 1'h0;
      write_enable_data_log_force[1879] <= 1'h0;
      write_enable_data_log_force[1880] <= 1'h0;
      write_enable_data_log_force[1881] <= 1'h0;
      write_enable_data_log_force[1882] <= 1'h0;
      write_enable_data_log_force[1883] <= 1'h0;
      write_enable_data_log_force[1884] <= 1'h0;
      write_enable_data_log_force[1885] <= 1'h0;
      write_enable_data_log_force[1886] <= 1'h0;
      write_enable_data_log_force[1887] <= 1'h0;
      write_enable_data_log_force[1888] <= 1'h0;
      write_enable_data_log_force[1889] <= 1'h0;
      write_enable_data_log_force[1890] <= 1'h0;
      write_enable_data_log_force[1891] <= 1'h0;
      write_enable_data_log_force[1892] <= 1'h0;
      write_enable_data_log_force[1893] <= 1'h0;
      write_enable_data_log_force[1894] <= 1'h0;
      write_enable_data_log_force[1895] <= 1'h0;
      write_enable_data_log_force[1896] <= 1'h0;
      write_enable_data_log_force[1897] <= 1'h0;
      write_enable_data_log_force[1898] <= 1'h0;
      write_enable_data_log_force[1899] <= 1'h0;
      write_enable_data_log_force[1900] <= 1'h0;
      write_enable_data_log_force[1901] <= 1'h0;
      write_enable_data_log_force[1902] <= 1'h0;
      write_enable_data_log_force[1903] <= 1'h0;
      write_enable_data_log_force[1904] <= 1'h0;
      write_enable_data_log_force[1905] <= 1'h0;
      write_enable_data_log_force[1906] <= 1'h0;
      write_enable_data_log_force[1907] <= 1'h0;
      write_enable_data_log_force[1908] <= 1'h0;
      write_enable_data_log_force[1909] <= 1'h0;
      write_enable_data_log_force[1910] <= 1'h0;
      write_enable_data_log_force[1911] <= 1'h0;
      write_enable_data_log_force[1912] <= 1'h0;
      write_enable_data_log_force[1913] <= 1'h0;
      write_enable_data_log_force[1914] <= 1'h0;
      write_enable_data_log_force[1915] <= 1'h0;
      write_enable_data_log_force[1916] <= 1'h0;
      write_enable_data_log_force[1917] <= 1'h0;
      write_enable_data_log_force[1918] <= 1'h0;
      write_enable_data_log_force[1919] <= 1'h0;
      write_enable_data_log_force[1920] <= 1'h0;
      write_enable_data_log_force[1921] <= 1'h0;
      write_enable_data_log_force[1922] <= 1'h0;
      write_enable_data_log_force[1923] <= 1'h0;
      write_enable_data_log_force[1924] <= 1'h0;
      write_enable_data_log_force[1925] <= 1'h0;
      write_enable_data_log_force[1926] <= 1'h0;
      write_enable_data_log_force[1927] <= 1'h0;
      write_enable_data_log_force[1928] <= 1'h0;
      write_enable_data_log_force[1929] <= 1'h0;
      write_enable_data_log_force[1930] <= 1'h0;
      write_enable_data_log_force[1931] <= 1'h0;
      write_enable_data_log_force[1932] <= 1'h0;
      write_enable_data_log_force[1933] <= 1'h0;
      write_enable_data_log_force[1934] <= 1'h0;
      write_enable_data_log_force[1935] <= 1'h0;
      write_enable_data_log_force[1936] <= 1'h0;
      write_enable_data_log_force[1937] <= 1'h0;
      write_enable_data_log_force[1938] <= 1'h0;
      write_enable_data_log_force[1939] <= 1'h0;
      write_enable_data_log_force[1940] <= 1'h0;
      write_enable_data_log_force[1941] <= 1'h0;
      write_enable_data_log_force[1942] <= 1'h0;
      write_enable_data_log_force[1943] <= 1'h0;
      write_enable_data_log_force[1944] <= 1'h0;
      write_enable_data_log_force[1945] <= 1'h0;
      write_enable_data_log_force[1946] <= 1'h0;
      write_enable_data_log_force[1947] <= 1'h0;
      write_enable_data_log_force[1948] <= 1'h0;
      write_enable_data_log_force[1949] <= 1'h0;
      write_enable_data_log_force[1950] <= 1'h0;
      write_enable_data_log_force[1951] <= 1'h0;
      write_enable_data_log_force[1952] <= 1'h0;
      write_enable_data_log_force[1953] <= 1'h0;
      write_enable_data_log_force[1954] <= 1'h0;
      write_enable_data_log_force[1955] <= 1'h0;
      write_enable_data_log_force[1956] <= 1'h0;
      write_enable_data_log_force[1957] <= 1'h0;
      write_enable_data_log_force[1958] <= 1'h0;
      write_enable_data_log_force[1959] <= 1'h0;
      write_enable_data_log_force[1960] <= 1'h0;
      write_enable_data_log_force[1961] <= 1'h0;
      write_enable_data_log_force[1962] <= 1'h0;
      write_enable_data_log_force[1963] <= 1'h0;
      write_enable_data_log_force[1964] <= 1'h0;
      write_enable_data_log_force[1965] <= 1'h0;
      write_enable_data_log_force[1966] <= 1'h0;
      write_enable_data_log_force[1967] <= 1'h0;
      write_enable_data_log_force[1968] <= 1'h0;
      write_enable_data_log_force[1969] <= 1'h0;
      write_enable_data_log_force[1970] <= 1'h0;
      write_enable_data_log_force[1971] <= 1'h0;
      write_enable_data_log_force[1972] <= 1'h0;
      write_enable_data_log_force[1973] <= 1'h0;
      write_enable_data_log_force[1974] <= 1'h0;
      write_enable_data_log_force[1975] <= 1'h0;
      write_enable_data_log_force[1976] <= 1'h0;
      write_enable_data_log_force[1977] <= 1'h0;
      write_enable_data_log_force[1978] <= 1'h0;
      write_enable_data_log_force[1979] <= 1'h0;
      write_enable_data_log_force[1980] <= 1'h0;
      write_enable_data_log_force[1981] <= 1'h0;
      write_enable_data_log_force[1982] <= 1'h0;
      write_enable_data_log_force[1983] <= 1'h0;
      write_enable_data_log_force[1984] <= 1'h0;
      write_enable_data_log_force[1985] <= 1'h0;
      write_enable_data_log_force[1986] <= 1'h0;
      write_enable_data_log_force[1987] <= 1'h0;
      write_enable_data_log_force[1988] <= 1'h0;
      write_enable_data_log_force[1989] <= 1'h0;
      write_enable_data_log_force[1990] <= 1'h0;
      write_enable_data_log_force[1991] <= 1'h0;
      write_enable_data_log_force[1992] <= 1'h0;
      write_enable_data_log_force[1993] <= 1'h0;
      write_enable_data_log_force[1994] <= 1'h0;
      write_enable_data_log_force[1995] <= 1'h0;
      write_enable_data_log_force[1996] <= 1'h0;
      write_enable_data_log_force[1997] <= 1'h0;
      write_enable_data_log_force[1998] <= 1'h0;
      write_enable_data_log_force[1999] <= 1'h0;
      write_enable_data_log_force[2000] <= 1'h0;
      write_enable_data_log_force[2001] <= 1'h0;
      write_enable_data_log_force[2002] <= 1'h0;
      write_enable_data_log_force[2003] <= 1'h0;
      write_enable_data_log_force[2004] <= 1'h0;
      write_enable_data_log_force[2005] <= 1'h0;
      write_enable_data_log_force[2006] <= 1'h0;
      write_enable_data_log_force[2007] <= 1'h0;
      write_enable_data_log_force[2008] <= 1'h0;
      write_enable_data_log_force[2009] <= 1'h0;
      write_enable_data_log_force[2010] <= 1'h0;
      write_enable_data_log_force[2011] <= 1'h0;
      write_enable_data_log_force[2012] <= 1'h0;
      write_enable_data_log_force[2013] <= 1'h0;
      write_enable_data_log_force[2014] <= 1'h0;
      write_enable_data_log_force[2015] <= 1'h0;
      write_enable_data_log_force[2016] <= 1'h0;
      write_enable_data_log_force[2017] <= 1'h0;
      write_enable_data_log_force[2018] <= 1'h0;
      write_enable_data_log_force[2019] <= 1'h0;
      write_enable_data_log_force[2020] <= 1'h0;
      write_enable_data_log_force[2021] <= 1'h0;
      write_enable_data_log_force[2022] <= 1'h0;
      write_enable_data_log_force[2023] <= 1'h0;
      write_enable_data_log_force[2024] <= 1'h0;
      write_enable_data_log_force[2025] <= 1'h0;
      write_enable_data_log_force[2026] <= 1'h0;
      write_enable_data_log_force[2027] <= 1'h0;
      write_enable_data_log_force[2028] <= 1'h0;
      write_enable_data_log_force[2029] <= 1'h0;
      write_enable_data_log_force[2030] <= 1'h0;
      write_enable_data_log_force[2031] <= 1'h0;
      write_enable_data_log_force[2032] <= 1'h0;
      write_enable_data_log_force[2033] <= 1'h0;
      write_enable_data_log_force[2034] <= 1'h0;
      write_enable_data_log_force[2035] <= 1'h0;
      write_enable_data_log_force[2036] <= 1'h0;
      write_enable_data_log_force[2037] <= 1'h0;
      write_enable_data_log_force[2038] <= 1'h0;
      write_enable_data_log_force[2039] <= 1'h0;
      write_enable_data_log_force[2040] <= 1'h0;
      write_enable_data_log_force[2041] <= 1'h0;
      write_enable_data_log_force[2042] <= 1'h0;
      write_enable_data_log_force[2043] <= 1'h0;
      write_enable_data_log_force[2044] <= 1'h0;
      write_enable_data_log_force[2045] <= 1'h0;
      write_enable_data_log_force[2046] <= 1'h0;
      write_enable_data_log_force[2047] <= 1'h0;
      write_enable_data_log_force[2048] <= 1'h0;
      write_enable_data_log_force[2049] <= 1'h0;
      write_enable_data_log_force[2050] <= 1'h0;
      write_enable_data_log_force[2051] <= 1'h0;
      write_enable_data_log_force[2052] <= 1'h0;
      write_enable_data_log_force[2053] <= 1'h0;
      write_enable_data_log_force[2054] <= 1'h0;
      write_enable_data_log_force[2055] <= 1'h0;
      write_enable_data_log_force[2056] <= 1'h0;
      write_enable_data_log_force[2057] <= 1'h0;
      write_enable_data_log_force[2058] <= 1'h0;
      write_enable_data_log_force[2059] <= 1'h0;
      write_enable_data_log_force[2060] <= 1'h0;
      write_enable_data_log_force[2061] <= 1'h0;
      write_enable_data_log_force[2062] <= 1'h0;
      write_enable_data_log_force[2063] <= 1'h0;
      write_enable_data_log_force[2064] <= 1'h0;
      write_enable_data_log_force[2065] <= 1'h0;
      write_enable_data_log_force[2066] <= 1'h0;
      write_enable_data_log_force[2067] <= 1'h0;
      write_enable_data_log_force[2068] <= 1'h0;
      write_enable_data_log_force[2069] <= 1'h0;
      write_enable_data_log_force[2070] <= 1'h0;
      write_enable_data_log_force[2071] <= 1'h0;
      write_enable_data_log_force[2072] <= 1'h0;
      write_enable_data_log_force[2073] <= 1'h0;
      write_enable_data_log_force[2074] <= 1'h0;
      write_enable_data_log_force[2075] <= 1'h0;
      write_enable_data_log_force[2076] <= 1'h0;
      write_enable_data_log_force[2077] <= 1'h0;
      write_enable_data_log_force[2078] <= 1'h0;
      write_enable_data_log_force[2079] <= 1'h0;
      write_enable_data_log_force[2080] <= 1'h0;
      write_enable_data_log_force[2081] <= 1'h0;
      write_enable_data_log_force[2082] <= 1'h0;
      write_enable_data_log_force[2083] <= 1'h0;
      write_enable_data_log_force[2084] <= 1'h0;
      write_enable_data_log_force[2085] <= 1'h0;
      write_enable_data_log_force[2086] <= 1'h0;
      write_enable_data_log_force[2087] <= 1'h0;
      write_enable_data_log_force[2088] <= 1'h0;
      write_enable_data_log_force[2089] <= 1'h0;
      write_enable_data_log_force[2090] <= 1'h0;
      write_enable_data_log_force[2091] <= 1'h0;
      write_enable_data_log_force[2092] <= 1'h0;
      write_enable_data_log_force[2093] <= 1'h0;
      write_enable_data_log_force[2094] <= 1'h0;
      write_enable_data_log_force[2095] <= 1'h0;
      write_enable_data_log_force[2096] <= 1'h0;
      write_enable_data_log_force[2097] <= 1'h0;
      write_enable_data_log_force[2098] <= 1'h0;
      write_enable_data_log_force[2099] <= 1'h0;
      write_enable_data_log_force[2100] <= 1'h0;
      write_enable_data_log_force[2101] <= 1'h0;
      write_enable_data_log_force[2102] <= 1'h0;
      write_enable_data_log_force[2103] <= 1'h0;
      write_enable_data_log_force[2104] <= 1'h0;
      write_enable_data_log_force[2105] <= 1'h0;
      write_enable_data_log_force[2106] <= 1'h0;
      write_enable_data_log_force[2107] <= 1'h0;
      write_enable_data_log_force[2108] <= 1'h0;
      write_enable_data_log_force[2109] <= 1'h0;
      write_enable_data_log_force[2110] <= 1'h0;
      write_enable_data_log_force[2111] <= 1'h0;
      write_enable_data_log_force[2112] <= 1'h0;
      write_enable_data_log_force[2113] <= 1'h0;
      write_enable_data_log_force[2114] <= 1'h0;
      write_enable_data_log_force[2115] <= 1'h0;
      write_enable_data_log_force[2116] <= 1'h0;
      write_enable_data_log_force[2117] <= 1'h0;
      write_enable_data_log_force[2118] <= 1'h0;
      write_enable_data_log_force[2119] <= 1'h0;
      write_enable_data_log_force[2120] <= 1'h0;
      write_enable_data_log_force[2121] <= 1'h0;
      write_enable_data_log_force[2122] <= 1'h0;
      write_enable_data_log_force[2123] <= 1'h0;
      write_enable_data_log_force[2124] <= 1'h0;
      write_enable_data_log_force[2125] <= 1'h0;
      write_enable_data_log_force[2126] <= 1'h0;
      write_enable_data_log_force[2127] <= 1'h0;
      write_enable_data_log_force[2128] <= 1'h0;
      write_enable_data_log_force[2129] <= 1'h0;
      write_enable_data_log_force[2130] <= 1'h0;
      write_enable_data_log_force[2131] <= 1'h0;
      write_enable_data_log_force[2132] <= 1'h0;
      write_enable_data_log_force[2133] <= 1'h0;
      write_enable_data_log_force[2134] <= 1'h0;
      write_enable_data_log_force[2135] <= 1'h0;
      write_enable_data_log_force[2136] <= 1'h0;
      write_enable_data_log_force[2137] <= 1'h0;
      write_enable_data_log_force[2138] <= 1'h0;
      write_enable_data_log_force[2139] <= 1'h0;
      write_enable_data_log_force[2140] <= 1'h0;
      write_enable_data_log_force[2141] <= 1'h0;
      write_enable_data_log_force[2142] <= 1'h0;
      write_enable_data_log_force[2143] <= 1'h0;
      write_enable_data_log_force[2144] <= 1'h0;
      write_enable_data_log_force[2145] <= 1'h0;
      write_enable_data_log_force[2146] <= 1'h0;
      write_enable_data_log_force[2147] <= 1'h0;
      write_enable_data_log_force[2148] <= 1'h0;
      write_enable_data_log_force[2149] <= 1'h0;
      write_enable_data_log_force[2150] <= 1'h0;
      write_enable_data_log_force[2151] <= 1'h0;
      write_enable_data_log_force[2152] <= 1'h0;
      write_enable_data_log_force[2153] <= 1'h0;
      write_enable_data_log_force[2154] <= 1'h0;
      write_enable_data_log_force[2155] <= 1'h0;
      write_enable_data_log_force[2156] <= 1'h0;
      write_enable_data_log_force[2157] <= 1'h0;
      write_enable_data_log_force[2158] <= 1'h0;
      write_enable_data_log_force[2159] <= 1'h0;
      write_enable_data_log_force[2160] <= 1'h0;
      write_enable_data_log_force[2161] <= 1'h0;
      write_enable_data_log_force[2162] <= 1'h0;
      write_enable_data_log_force[2163] <= 1'h0;
      write_enable_data_log_force[2164] <= 1'h0;
      write_enable_data_log_force[2165] <= 1'h0;
      write_enable_data_log_force[2166] <= 1'h0;
      write_enable_data_log_force[2167] <= 1'h0;
      write_enable_data_log_force[2168] <= 1'h0;
      write_enable_data_log_force[2169] <= 1'h0;
      write_enable_data_log_force[2170] <= 1'h0;
      write_enable_data_log_force[2171] <= 1'h0;
      write_enable_data_log_force[2172] <= 1'h0;
      write_enable_data_log_force[2173] <= 1'h0;
      write_enable_data_log_force[2174] <= 1'h0;
      write_enable_data_log_force[2175] <= 1'h0;
      write_enable_data_log_force[2176] <= 1'h0;
      write_enable_data_log_force[2177] <= 1'h0;
      write_enable_data_log_force[2178] <= 1'h0;
      write_enable_data_log_force[2179] <= 1'h0;
      write_enable_data_log_force[2180] <= 1'h0;
      write_enable_data_log_force[2181] <= 1'h0;
      write_enable_data_log_force[2182] <= 1'h0;
      write_enable_data_log_force[2183] <= 1'h0;
      write_enable_data_log_force[2184] <= 1'h0;
      write_enable_data_log_force[2185] <= 1'h0;
      write_enable_data_log_force[2186] <= 1'h0;
      write_enable_data_log_force[2187] <= 1'h0;
      write_enable_data_log_force[2188] <= 1'h0;
      write_enable_data_log_force[2189] <= 1'h0;
      write_enable_data_log_force[2190] <= 1'h0;
      write_enable_data_log_force[2191] <= 1'h0;
      write_enable_data_log_force[2192] <= 1'h0;
      write_enable_data_log_force[2193] <= 1'h0;
      write_enable_data_log_force[2194] <= 1'h0;
      write_enable_data_log_force[2195] <= 1'h0;
      write_enable_data_log_force[2196] <= 1'h0;
      write_enable_data_log_force[2197] <= 1'h0;
      write_enable_data_log_force[2198] <= 1'h0;
      write_enable_data_log_force[2199] <= 1'h0;
      write_enable_data_log_force[2200] <= 1'h0;
      write_enable_data_log_force[2201] <= 1'h0;
      write_enable_data_log_force[2202] <= 1'h0;
      write_enable_data_log_force[2203] <= 1'h0;
      write_enable_data_log_force[2204] <= 1'h0;
      write_enable_data_log_force[2205] <= 1'h0;
      write_enable_data_log_force[2206] <= 1'h0;
      write_enable_data_log_force[2207] <= 1'h0;
      write_enable_data_log_force[2208] <= 1'h0;
      write_enable_data_log_force[2209] <= 1'h0;
      write_enable_data_log_force[2210] <= 1'h0;
      write_enable_data_log_force[2211] <= 1'h0;
      write_enable_data_log_force[2212] <= 1'h0;
      write_enable_data_log_force[2213] <= 1'h0;
      write_enable_data_log_force[2214] <= 1'h0;
      write_enable_data_log_force[2215] <= 1'h0;
      write_enable_data_log_force[2216] <= 1'h0;
      write_enable_data_log_force[2217] <= 1'h0;
      write_enable_data_log_force[2218] <= 1'h0;
      write_enable_data_log_force[2219] <= 1'h0;
      write_enable_data_log_force[2220] <= 1'h0;
      write_enable_data_log_force[2221] <= 1'h0;
      write_enable_data_log_force[2222] <= 1'h0;
      write_enable_data_log_force[2223] <= 1'h0;
      write_enable_data_log_force[2224] <= 1'h0;
      write_enable_data_log_force[2225] <= 1'h0;
      write_enable_data_log_force[2226] <= 1'h0;
      write_enable_data_log_force[2227] <= 1'h0;
      write_enable_data_log_force[2228] <= 1'h0;
      write_enable_data_log_force[2229] <= 1'h0;
      write_enable_data_log_force[2230] <= 1'h0;
      write_enable_data_log_force[2231] <= 1'h0;
      write_enable_data_log_force[2232] <= 1'h0;
      write_enable_data_log_force[2233] <= 1'h0;
      write_enable_data_log_force[2234] <= 1'h0;
      write_enable_data_log_force[2235] <= 1'h0;
      write_enable_data_log_force[2236] <= 1'h0;
      write_enable_data_log_force[2237] <= 1'h0;
      write_enable_data_log_force[2238] <= 1'h0;
      write_enable_data_log_force[2239] <= 1'h0;
      write_enable_data_log_force[2240] <= 1'h0;
      write_enable_data_log_force[2241] <= 1'h0;
      write_enable_data_log_force[2242] <= 1'h0;
      write_enable_data_log_force[2243] <= 1'h0;
      write_enable_data_log_force[2244] <= 1'h0;
      write_enable_data_log_force[2245] <= 1'h0;
      write_enable_data_log_force[2246] <= 1'h0;
      write_enable_data_log_force[2247] <= 1'h0;
      write_enable_data_log_force[2248] <= 1'h0;
      write_enable_data_log_force[2249] <= 1'h0;
      write_enable_data_log_force[2250] <= 1'h0;
      write_enable_data_log_force[2251] <= 1'h0;
      write_enable_data_log_force[2252] <= 1'h0;
      write_enable_data_log_force[2253] <= 1'h0;
      write_enable_data_log_force[2254] <= 1'h0;
      write_enable_data_log_force[2255] <= 1'h0;
      write_enable_data_log_force[2256] <= 1'h0;
      write_enable_data_log_force[2257] <= 1'h0;
      write_enable_data_log_force[2258] <= 1'h0;
      write_enable_data_log_force[2259] <= 1'h0;
      write_enable_data_log_force[2260] <= 1'h0;
      write_enable_data_log_force[2261] <= 1'h0;
      write_enable_data_log_force[2262] <= 1'h0;
      write_enable_data_log_force[2263] <= 1'h0;
      write_enable_data_log_force[2264] <= 1'h0;
      write_enable_data_log_force[2265] <= 1'h0;
      write_enable_data_log_force[2266] <= 1'h0;
      write_enable_data_log_force[2267] <= 1'h0;
      write_enable_data_log_force[2268] <= 1'h0;
      write_enable_data_log_force[2269] <= 1'h0;
      write_enable_data_log_force[2270] <= 1'h0;
      write_enable_data_log_force[2271] <= 1'h0;
      write_enable_data_log_force[2272] <= 1'h0;
      write_enable_data_log_force[2273] <= 1'h0;
      write_enable_data_log_force[2274] <= 1'h0;
      write_enable_data_log_force[2275] <= 1'h0;
      write_enable_data_log_force[2276] <= 1'h0;
      write_enable_data_log_force[2277] <= 1'h0;
      write_enable_data_log_force[2278] <= 1'h0;
      write_enable_data_log_force[2279] <= 1'h0;
      write_enable_data_log_force[2280] <= 1'h0;
      write_enable_data_log_force[2281] <= 1'h0;
      write_enable_data_log_force[2282] <= 1'h0;
      write_enable_data_log_force[2283] <= 1'h0;
      write_enable_data_log_force[2284] <= 1'h0;
      write_enable_data_log_force[2285] <= 1'h0;
      write_enable_data_log_force[2286] <= 1'h0;
      write_enable_data_log_force[2287] <= 1'h0;
      write_enable_data_log_force[2288] <= 1'h0;
      write_enable_data_log_force[2289] <= 1'h0;
      write_enable_data_log_force[2290] <= 1'h0;
      write_enable_data_log_force[2291] <= 1'h0;
      write_enable_data_log_force[2292] <= 1'h0;
      write_enable_data_log_force[2293] <= 1'h0;
      write_enable_data_log_force[2294] <= 1'h0;
      write_enable_data_log_force[2295] <= 1'h0;
      write_enable_data_log_force[2296] <= 1'h0;
      write_enable_data_log_force[2297] <= 1'h0;
      write_enable_data_log_force[2298] <= 1'h0;
      write_enable_data_log_force[2299] <= 1'h0;
      write_enable_data_log_force[2300] <= 1'h0;
      write_enable_data_log_force[2301] <= 1'h0;
      write_enable_data_log_force[2302] <= 1'h0;
      write_enable_data_log_force[2303] <= 1'h0;
      write_enable_data_log_force[2304] <= 1'h0;
      write_enable_data_log_force[2305] <= 1'h0;
      write_enable_data_log_force[2306] <= 1'h0;
      write_enable_data_log_force[2307] <= 1'h0;
      write_enable_data_log_force[2308] <= 1'h0;
      write_enable_data_log_force[2309] <= 1'h0;
      write_enable_data_log_force[2310] <= 1'h0;
      write_enable_data_log_force[2311] <= 1'h0;
      write_enable_data_log_force[2312] <= 1'h0;
      write_enable_data_log_force[2313] <= 1'h0;
      write_enable_data_log_force[2314] <= 1'h0;
      write_enable_data_log_force[2315] <= 1'h0;
      write_enable_data_log_force[2316] <= 1'h0;
      write_enable_data_log_force[2317] <= 1'h0;
      write_enable_data_log_force[2318] <= 1'h0;
      write_enable_data_log_force[2319] <= 1'h0;
      write_enable_data_log_force[2320] <= 1'h0;
      write_enable_data_log_force[2321] <= 1'h0;
      write_enable_data_log_force[2322] <= 1'h0;
      write_enable_data_log_force[2323] <= 1'h0;
      write_enable_data_log_force[2324] <= 1'h0;
      write_enable_data_log_force[2325] <= 1'h0;
      write_enable_data_log_force[2326] <= 1'h0;
      write_enable_data_log_force[2327] <= 1'h0;
      write_enable_data_log_force[2328] <= 1'h0;
      write_enable_data_log_force[2329] <= 1'h0;
      write_enable_data_log_force[2330] <= 1'h0;
      write_enable_data_log_force[2331] <= 1'h0;
      write_enable_data_log_force[2332] <= 1'h0;
      write_enable_data_log_force[2333] <= 1'h0;
      write_enable_data_log_force[2334] <= 1'h0;
      write_enable_data_log_force[2335] <= 1'h0;
      write_enable_data_log_force[2336] <= 1'h0;
      write_enable_data_log_force[2337] <= 1'h0;
      write_enable_data_log_force[2338] <= 1'h0;
      write_enable_data_log_force[2339] <= 1'h0;
      write_enable_data_log_force[2340] <= 1'h0;
      write_enable_data_log_force[2341] <= 1'h0;
      write_enable_data_log_force[2342] <= 1'h0;
      write_enable_data_log_force[2343] <= 1'h0;
      write_enable_data_log_force[2344] <= 1'h0;
      write_enable_data_log_force[2345] <= 1'h0;
      write_enable_data_log_force[2346] <= 1'h0;
      write_enable_data_log_force[2347] <= 1'h0;
      write_enable_data_log_force[2348] <= 1'h0;
      write_enable_data_log_force[2349] <= 1'h0;
      write_enable_data_log_force[2350] <= 1'h0;
      write_enable_data_log_force[2351] <= 1'h0;
      write_enable_data_log_force[2352] <= 1'h0;
      write_enable_data_log_force[2353] <= 1'h0;
      write_enable_data_log_force[2354] <= 1'h0;
      write_enable_data_log_force[2355] <= 1'h0;
      write_enable_data_log_force[2356] <= 1'h0;
      write_enable_data_log_force[2357] <= 1'h0;
      write_enable_data_log_force[2358] <= 1'h0;
      write_enable_data_log_force[2359] <= 1'h0;
      write_enable_data_log_force[2360] <= 1'h0;
      write_enable_data_log_force[2361] <= 1'h0;
      write_enable_data_log_force[2362] <= 1'h0;
      write_enable_data_log_force[2363] <= 1'h0;
      write_enable_data_log_force[2364] <= 1'h0;
      write_enable_data_log_force[2365] <= 1'h0;
      write_enable_data_log_force[2366] <= 1'h0;
      write_enable_data_log_force[2367] <= 1'h0;
      write_enable_data_log_force[2368] <= 1'h0;
      write_enable_data_log_force[2369] <= 1'h0;
      write_enable_data_log_force[2370] <= 1'h0;
      write_enable_data_log_force[2371] <= 1'h0;
      write_enable_data_log_force[2372] <= 1'h0;
      write_enable_data_log_force[2373] <= 1'h0;
      write_enable_data_log_force[2374] <= 1'h0;
      write_enable_data_log_force[2375] <= 1'h0;
      write_enable_data_log_force[2376] <= 1'h0;
      write_enable_data_log_force[2377] <= 1'h0;
      write_enable_data_log_force[2378] <= 1'h0;
      write_enable_data_log_force[2379] <= 1'h0;
      write_enable_data_log_force[2380] <= 1'h0;
      write_enable_data_log_force[2381] <= 1'h0;
      write_enable_data_log_force[2382] <= 1'h0;
      write_enable_data_log_force[2383] <= 1'h0;
      write_enable_data_log_force[2384] <= 1'h0;
      write_enable_data_log_force[2385] <= 1'h0;
      write_enable_data_log_force[2386] <= 1'h0;
      write_enable_data_log_force[2387] <= 1'h0;
      write_enable_data_log_force[2388] <= 1'h0;
      write_enable_data_log_force[2389] <= 1'h0;
      write_enable_data_log_force[2390] <= 1'h0;
      write_enable_data_log_force[2391] <= 1'h0;
      write_enable_data_log_force[2392] <= 1'h0;
      write_enable_data_log_force[2393] <= 1'h0;
      write_enable_data_log_force[2394] <= 1'h0;
      write_enable_data_log_force[2395] <= 1'h0;
      write_enable_data_log_force[2396] <= 1'h0;
      write_enable_data_log_force[2397] <= 1'h0;
      write_enable_data_log_force[2398] <= 1'h0;
      write_enable_data_log_force[2399] <= 1'h0;
      write_enable_data_log_force[2400] <= 1'h0;
      write_enable_data_log_force[2401] <= 1'h0;
      write_enable_data_log_force[2402] <= 1'h0;
      write_enable_data_log_force[2403] <= 1'h0;
      write_enable_data_log_force[2404] <= 1'h0;
      write_enable_data_log_force[2405] <= 1'h0;
      write_enable_data_log_force[2406] <= 1'h0;
      write_enable_data_log_force[2407] <= 1'h0;
      write_enable_data_log_force[2408] <= 1'h0;
      write_enable_data_log_force[2409] <= 1'h0;
      write_enable_data_log_force[2410] <= 1'h0;
      write_enable_data_log_force[2411] <= 1'h0;
      write_enable_data_log_force[2412] <= 1'h0;
      write_enable_data_log_force[2413] <= 1'h0;
      write_enable_data_log_force[2414] <= 1'h0;
      write_enable_data_log_force[2415] <= 1'h0;
      write_enable_data_log_force[2416] <= 1'h0;
      write_enable_data_log_force[2417] <= 1'h0;
      write_enable_data_log_force[2418] <= 1'h0;
      write_enable_data_log_force[2419] <= 1'h0;
      write_enable_data_log_force[2420] <= 1'h0;
      write_enable_data_log_force[2421] <= 1'h0;
      write_enable_data_log_force[2422] <= 1'h0;
      write_enable_data_log_force[2423] <= 1'h0;
      write_enable_data_log_force[2424] <= 1'h0;
      write_enable_data_log_force[2425] <= 1'h0;
      write_enable_data_log_force[2426] <= 1'h0;
      write_enable_data_log_force[2427] <= 1'h0;
      write_enable_data_log_force[2428] <= 1'h0;
      write_enable_data_log_force[2429] <= 1'h0;
      write_enable_data_log_force[2430] <= 1'h0;
      write_enable_data_log_force[2431] <= 1'h0;
      write_enable_data_log_force[2432] <= 1'h0;
      write_enable_data_log_force[2433] <= 1'h0;
      write_enable_data_log_force[2434] <= 1'h0;
      write_enable_data_log_force[2435] <= 1'h0;
      write_enable_data_log_force[2436] <= 1'h0;
      write_enable_data_log_force[2437] <= 1'h0;
      write_enable_data_log_force[2438] <= 1'h0;
      write_enable_data_log_force[2439] <= 1'h0;
      write_enable_data_log_force[2440] <= 1'h0;
      write_enable_data_log_force[2441] <= 1'h0;
      write_enable_data_log_force[2442] <= 1'h0;
      write_enable_data_log_force[2443] <= 1'h0;
      write_enable_data_log_force[2444] <= 1'h0;
      write_enable_data_log_force[2445] <= 1'h0;
      write_enable_data_log_force[2446] <= 1'h0;
      write_enable_data_log_force[2447] <= 1'h0;
      write_enable_data_log_force[2448] <= 1'h0;
      write_enable_data_log_force[2449] <= 1'h0;
      write_enable_data_log_force[2450] <= 1'h0;
      write_enable_data_log_force[2451] <= 1'h0;
      write_enable_data_log_force[2452] <= 1'h0;
      write_enable_data_log_force[2453] <= 1'h0;
      write_enable_data_log_force[2454] <= 1'h0;
      write_enable_data_log_force[2455] <= 1'h0;
      write_enable_data_log_force[2456] <= 1'h0;
      write_enable_data_log_force[2457] <= 1'h0;
      write_enable_data_log_force[2458] <= 1'h0;
      write_enable_data_log_force[2459] <= 1'h0;
      write_enable_data_log_force[2460] <= 1'h0;
      write_enable_data_log_force[2461] <= 1'h0;
      write_enable_data_log_force[2462] <= 1'h0;
      write_enable_data_log_force[2463] <= 1'h0;
      write_enable_data_log_force[2464] <= 1'h0;
      write_enable_data_log_force[2465] <= 1'h0;
      write_enable_data_log_force[2466] <= 1'h0;
      write_enable_data_log_force[2467] <= 1'h0;
      write_enable_data_log_force[2468] <= 1'h0;
      write_enable_data_log_force[2469] <= 1'h0;
      write_enable_data_log_force[2470] <= 1'h0;
      write_enable_data_log_force[2471] <= 1'h0;
      write_enable_data_log_force[2472] <= 1'h0;
      write_enable_data_log_force[2473] <= 1'h0;
      write_enable_data_log_force[2474] <= 1'h0;
      write_enable_data_log_force[2475] <= 1'h0;
      write_enable_data_log_force[2476] <= 1'h0;
      write_enable_data_log_force[2477] <= 1'h0;
      write_enable_data_log_force[2478] <= 1'h0;
      write_enable_data_log_force[2479] <= 1'h0;
      write_enable_data_log_force[2480] <= 1'h0;
      write_enable_data_log_force[2481] <= 1'h0;
      write_enable_data_log_force[2482] <= 1'h0;
      write_enable_data_log_force[2483] <= 1'h0;
      write_enable_data_log_force[2484] <= 1'h0;
      write_enable_data_log_force[2485] <= 1'h0;
      write_enable_data_log_force[2486] <= 1'h0;
      write_enable_data_log_force[2487] <= 1'h0;
      write_enable_data_log_force[2488] <= 1'h0;
      write_enable_data_log_force[2489] <= 1'h0;
      write_enable_data_log_force[2490] <= 1'h0;
      write_enable_data_log_force[2491] <= 1'h0;
      write_enable_data_log_force[2492] <= 1'h0;
      write_enable_data_log_force[2493] <= 1'h0;
      write_enable_data_log_force[2494] <= 1'h0;
      write_enable_data_log_force[2495] <= 1'h0;
      write_enable_data_log_force[2496] <= 1'h0;
      write_enable_data_log_force[2497] <= 1'h0;
      write_enable_data_log_force[2498] <= 1'h0;
      write_enable_data_log_force[2499] <= 1'h0;
      write_enable_data_log_force[2500] <= 1'h0;
      write_enable_data_log_force[2501] <= 1'h0;
      write_enable_data_log_force[2502] <= 1'h0;
      write_enable_data_log_force[2503] <= 1'h0;
      write_enable_data_log_force[2504] <= 1'h0;
      write_enable_data_log_force[2505] <= 1'h0;
      write_enable_data_log_force[2506] <= 1'h0;
      write_enable_data_log_force[2507] <= 1'h0;
      write_enable_data_log_force[2508] <= 1'h0;
      write_enable_data_log_force[2509] <= 1'h0;
      write_enable_data_log_force[2510] <= 1'h0;
      write_enable_data_log_force[2511] <= 1'h0;
      write_enable_data_log_force[2512] <= 1'h0;
      write_enable_data_log_force[2513] <= 1'h0;
      write_enable_data_log_force[2514] <= 1'h0;
      write_enable_data_log_force[2515] <= 1'h0;
      write_enable_data_log_force[2516] <= 1'h0;
      write_enable_data_log_force[2517] <= 1'h0;
      write_enable_data_log_force[2518] <= 1'h0;
      write_enable_data_log_force[2519] <= 1'h0;
      write_enable_data_log_force[2520] <= 1'h0;
      write_enable_data_log_force[2521] <= 1'h0;
      write_enable_data_log_force[2522] <= 1'h0;
      write_enable_data_log_force[2523] <= 1'h0;
      write_enable_data_log_force[2524] <= 1'h0;
      write_enable_data_log_force[2525] <= 1'h0;
      write_enable_data_log_force[2526] <= 1'h0;
      write_enable_data_log_force[2527] <= 1'h0;
      write_enable_data_log_force[2528] <= 1'h0;
      write_enable_data_log_force[2529] <= 1'h0;
      write_enable_data_log_force[2530] <= 1'h0;
      write_enable_data_log_force[2531] <= 1'h0;
      write_enable_data_log_force[2532] <= 1'h0;
      write_enable_data_log_force[2533] <= 1'h0;
      write_enable_data_log_force[2534] <= 1'h0;
      write_enable_data_log_force[2535] <= 1'h0;
      write_enable_data_log_force[2536] <= 1'h0;
      write_enable_data_log_force[2537] <= 1'h0;
      write_enable_data_log_force[2538] <= 1'h0;
      write_enable_data_log_force[2539] <= 1'h0;
      write_enable_data_log_force[2540] <= 1'h0;
      write_enable_data_log_force[2541] <= 1'h0;
      write_enable_data_log_force[2542] <= 1'h0;
      write_enable_data_log_force[2543] <= 1'h0;
      write_enable_data_log_force[2544] <= 1'h0;
      write_enable_data_log_force[2545] <= 1'h0;
      write_enable_data_log_force[2546] <= 1'h0;
      write_enable_data_log_force[2547] <= 1'h0;
      write_enable_data_log_force[2548] <= 1'h0;
      write_enable_data_log_force[2549] <= 1'h0;
      write_enable_data_log_force[2550] <= 1'h0;
      write_enable_data_log_force[2551] <= 1'h0;
      write_enable_data_log_force[2552] <= 1'h0;
      write_enable_data_log_force[2553] <= 1'h0;
      write_enable_data_log_force[2554] <= 1'h0;
      write_enable_data_log_force[2555] <= 1'h0;
      write_enable_data_log_force[2556] <= 1'h0;
      write_enable_data_log_force[2557] <= 1'h0;
      write_enable_data_log_force[2558] <= 1'h0;
      write_enable_data_log_force[2559] <= 1'h0;
      write_enable_data_log_force[2560] <= 1'h0;
      write_enable_data_log_force[2561] <= 1'h0;
      write_enable_data_log_force[2562] <= 1'h0;
      write_enable_data_log_force[2563] <= 1'h0;
      write_enable_data_log_force[2564] <= 1'h0;
      write_enable_data_log_force[2565] <= 1'h0;
      write_enable_data_log_force[2566] <= 1'h0;
      write_enable_data_log_force[2567] <= 1'h0;
      write_enable_data_log_force[2568] <= 1'h0;
      write_enable_data_log_force[2569] <= 1'h0;
      write_enable_data_log_force[2570] <= 1'h0;
      write_enable_data_log_force[2571] <= 1'h0;
      write_enable_data_log_force[2572] <= 1'h0;
      write_enable_data_log_force[2573] <= 1'h0;
      write_enable_data_log_force[2574] <= 1'h0;
      write_enable_data_log_force[2575] <= 1'h0;
      write_enable_data_log_force[2576] <= 1'h0;
      write_enable_data_log_force[2577] <= 1'h0;
      write_enable_data_log_force[2578] <= 1'h0;
      write_enable_data_log_force[2579] <= 1'h0;
      write_enable_data_log_force[2580] <= 1'h0;
      write_enable_data_log_force[2581] <= 1'h0;
      write_enable_data_log_force[2582] <= 1'h0;
      write_enable_data_log_force[2583] <= 1'h0;
      write_enable_data_log_force[2584] <= 1'h0;
      write_enable_data_log_force[2585] <= 1'h0;
      write_enable_data_log_force[2586] <= 1'h0;
      write_enable_data_log_force[2587] <= 1'h0;
      write_enable_data_log_force[2588] <= 1'h0;
      write_enable_data_log_force[2589] <= 1'h0;
      write_enable_data_log_force[2590] <= 1'h0;
      write_enable_data_log_force[2591] <= 1'h0;
      write_enable_data_log_force[2592] <= 1'h0;
      write_enable_data_log_force[2593] <= 1'h0;
      write_enable_data_log_force[2594] <= 1'h0;
      write_enable_data_log_force[2595] <= 1'h0;
      write_enable_data_log_force[2596] <= 1'h0;
      write_enable_data_log_force[2597] <= 1'h0;
      write_enable_data_log_force[2598] <= 1'h0;
      write_enable_data_log_force[2599] <= 1'h0;
      write_enable_data_log_force[2600] <= 1'h0;
      write_enable_data_log_force[2601] <= 1'h0;
      write_enable_data_log_force[2602] <= 1'h0;
      write_enable_data_log_force[2603] <= 1'h0;
      write_enable_data_log_force[2604] <= 1'h0;
      write_enable_data_log_force[2605] <= 1'h0;
      write_enable_data_log_force[2606] <= 1'h0;
      write_enable_data_log_force[2607] <= 1'h0;
      write_enable_data_log_force[2608] <= 1'h0;
      write_enable_data_log_force[2609] <= 1'h0;
      write_enable_data_log_force[2610] <= 1'h0;
      write_enable_data_log_force[2611] <= 1'h0;
      write_enable_data_log_force[2612] <= 1'h0;
      write_enable_data_log_force[2613] <= 1'h0;
      write_enable_data_log_force[2614] <= 1'h0;
      write_enable_data_log_force[2615] <= 1'h0;
      write_enable_data_log_force[2616] <= 1'h0;
      write_enable_data_log_force[2617] <= 1'h0;
      write_enable_data_log_force[2618] <= 1'h0;
      write_enable_data_log_force[2619] <= 1'h0;
      write_enable_data_log_force[2620] <= 1'h0;
      write_enable_data_log_force[2621] <= 1'h0;
      write_enable_data_log_force[2622] <= 1'h0;
      write_enable_data_log_force[2623] <= 1'h0;
      write_enable_data_log_force[2624] <= 1'h0;
      write_enable_data_log_force[2625] <= 1'h0;
      write_enable_data_log_force[2626] <= 1'h0;
      write_enable_data_log_force[2627] <= 1'h0;
      write_enable_data_log_force[2628] <= 1'h0;
      write_enable_data_log_force[2629] <= 1'h0;
      write_enable_data_log_force[2630] <= 1'h0;
      write_enable_data_log_force[2631] <= 1'h0;
      write_enable_data_log_force[2632] <= 1'h0;
      write_enable_data_log_force[2633] <= 1'h0;
      write_enable_data_log_force[2634] <= 1'h0;
      write_enable_data_log_force[2635] <= 1'h0;
      write_enable_data_log_force[2636] <= 1'h0;
      write_enable_data_log_force[2637] <= 1'h0;
      write_enable_data_log_force[2638] <= 1'h0;
      write_enable_data_log_force[2639] <= 1'h0;
      write_enable_data_log_force[2640] <= 1'h0;
      write_enable_data_log_force[2641] <= 1'h0;
      write_enable_data_log_force[2642] <= 1'h0;
      write_enable_data_log_force[2643] <= 1'h0;
      write_enable_data_log_force[2644] <= 1'h0;
      write_enable_data_log_force[2645] <= 1'h0;
      write_enable_data_log_force[2646] <= 1'h0;
      write_enable_data_log_force[2647] <= 1'h0;
      write_enable_data_log_force[2648] <= 1'h0;
      write_enable_data_log_force[2649] <= 1'h0;
      write_enable_data_log_force[2650] <= 1'h0;
      write_enable_data_log_force[2651] <= 1'h0;
      write_enable_data_log_force[2652] <= 1'h0;
      write_enable_data_log_force[2653] <= 1'h0;
      write_enable_data_log_force[2654] <= 1'h0;
      write_enable_data_log_force[2655] <= 1'h0;
      write_enable_data_log_force[2656] <= 1'h0;
      write_enable_data_log_force[2657] <= 1'h0;
      write_enable_data_log_force[2658] <= 1'h0;
      write_enable_data_log_force[2659] <= 1'h0;
      write_enable_data_log_force[2660] <= 1'h0;
      write_enable_data_log_force[2661] <= 1'h0;
      write_enable_data_log_force[2662] <= 1'h0;
      write_enable_data_log_force[2663] <= 1'h0;
      write_enable_data_log_force[2664] <= 1'h0;
      write_enable_data_log_force[2665] <= 1'h0;
      write_enable_data_log_force[2666] <= 1'h0;
      write_enable_data_log_force[2667] <= 1'h0;
      write_enable_data_log_force[2668] <= 1'h0;
      write_enable_data_log_force[2669] <= 1'h0;
      write_enable_data_log_force[2670] <= 1'h0;
      write_enable_data_log_force[2671] <= 1'h0;
      write_enable_data_log_force[2672] <= 1'h0;
      write_enable_data_log_force[2673] <= 1'h0;
      write_enable_data_log_force[2674] <= 1'h0;
      write_enable_data_log_force[2675] <= 1'h0;
      write_enable_data_log_force[2676] <= 1'h0;
      write_enable_data_log_force[2677] <= 1'h0;
      write_enable_data_log_force[2678] <= 1'h0;
      write_enable_data_log_force[2679] <= 1'h0;
      write_enable_data_log_force[2680] <= 1'h0;
      write_enable_data_log_force[2681] <= 1'h0;
      write_enable_data_log_force[2682] <= 1'h0;
      write_enable_data_log_force[2683] <= 1'h0;
      write_enable_data_log_force[2684] <= 1'h0;
      write_enable_data_log_force[2685] <= 1'h0;
      write_enable_data_log_force[2686] <= 1'h0;
      write_enable_data_log_force[2687] <= 1'h0;
      write_enable_data_log_force[2688] <= 1'h0;
      write_enable_data_log_force[2689] <= 1'h0;
      write_enable_data_log_force[2690] <= 1'h0;
      write_enable_data_log_force[2691] <= 1'h0;
      write_enable_data_log_force[2692] <= 1'h0;
      write_enable_data_log_force[2693] <= 1'h0;
      write_enable_data_log_force[2694] <= 1'h0;
      write_enable_data_log_force[2695] <= 1'h0;
      write_enable_data_log_force[2696] <= 1'h0;
      write_enable_data_log_force[2697] <= 1'h0;
      write_enable_data_log_force[2698] <= 1'h0;
      write_enable_data_log_force[2699] <= 1'h0;
      write_enable_data_log_force[2700] <= 1'h0;
      write_enable_data_log_force[2701] <= 1'h0;
      write_enable_data_log_force[2702] <= 1'h0;
      write_enable_data_log_force[2703] <= 1'h0;
      write_enable_data_log_force[2704] <= 1'h0;
      write_enable_data_log_force[2705] <= 1'h0;
      write_enable_data_log_force[2706] <= 1'h0;
      write_enable_data_log_force[2707] <= 1'h0;
      write_enable_data_log_force[2708] <= 1'h0;
      write_enable_data_log_force[2709] <= 1'h0;
      write_enable_data_log_force[2710] <= 1'h0;
      write_enable_data_log_force[2711] <= 1'h0;
      write_enable_data_log_force[2712] <= 1'h0;
      write_enable_data_log_force[2713] <= 1'h0;
      write_enable_data_log_force[2714] <= 1'h0;
      write_enable_data_log_force[2715] <= 1'h0;
      write_enable_data_log_force[2716] <= 1'h0;
      write_enable_data_log_force[2717] <= 1'h0;
      write_enable_data_log_force[2718] <= 1'h0;
      write_enable_data_log_force[2719] <= 1'h0;
      write_enable_data_log_force[2720] <= 1'h0;
      write_enable_data_log_force[2721] <= 1'h0;
      write_enable_data_log_force[2722] <= 1'h0;
      write_enable_data_log_force[2723] <= 1'h0;
      write_enable_data_log_force[2724] <= 1'h0;
      write_enable_data_log_force[2725] <= 1'h0;
      write_enable_data_log_force[2726] <= 1'h0;
      write_enable_data_log_force[2727] <= 1'h0;
      write_enable_data_log_force[2728] <= 1'h0;
      write_enable_data_log_force[2729] <= 1'h0;
      write_enable_data_log_force[2730] <= 1'h0;
      write_enable_data_log_force[2731] <= 1'h0;
      write_enable_data_log_force[2732] <= 1'h0;
      write_enable_data_log_force[2733] <= 1'h0;
      write_enable_data_log_force[2734] <= 1'h0;
      write_enable_data_log_force[2735] <= 1'h0;
      write_enable_data_log_force[2736] <= 1'h0;
      write_enable_data_log_force[2737] <= 1'h0;
      write_enable_data_log_force[2738] <= 1'h0;
      write_enable_data_log_force[2739] <= 1'h0;
      write_enable_data_log_force[2740] <= 1'h0;
      write_enable_data_log_force[2741] <= 1'h0;
      write_enable_data_log_force[2742] <= 1'h0;
      write_enable_data_log_force[2743] <= 1'h0;
      write_enable_data_log_force[2744] <= 1'h0;
      write_enable_data_log_force[2745] <= 1'h0;
      write_enable_data_log_force[2746] <= 1'h0;
      write_enable_data_log_force[2747] <= 1'h0;
      write_enable_data_log_force[2748] <= 1'h0;
      write_enable_data_log_force[2749] <= 1'h0;
      write_enable_data_log_force[2750] <= 1'h0;
      write_enable_data_log_force[2751] <= 1'h0;
      write_enable_data_log_force[2752] <= 1'h0;
      write_enable_data_log_force[2753] <= 1'h0;
      write_enable_data_log_force[2754] <= 1'h0;
      write_enable_data_log_force[2755] <= 1'h0;
      write_enable_data_log_force[2756] <= 1'h0;
      write_enable_data_log_force[2757] <= 1'h0;
      write_enable_data_log_force[2758] <= 1'h0;
      write_enable_data_log_force[2759] <= 1'h0;
      write_enable_data_log_force[2760] <= 1'h0;
      write_enable_data_log_force[2761] <= 1'h0;
      write_enable_data_log_force[2762] <= 1'h0;
      write_enable_data_log_force[2763] <= 1'h0;
      write_enable_data_log_force[2764] <= 1'h0;
      write_enable_data_log_force[2765] <= 1'h0;
      write_enable_data_log_force[2766] <= 1'h0;
      write_enable_data_log_force[2767] <= 1'h0;
      write_enable_data_log_force[2768] <= 1'h0;
      write_enable_data_log_force[2769] <= 1'h0;
      write_enable_data_log_force[2770] <= 1'h0;
      write_enable_data_log_force[2771] <= 1'h0;
      write_enable_data_log_force[2772] <= 1'h0;
      write_enable_data_log_force[2773] <= 1'h0;
      write_enable_data_log_force[2774] <= 1'h0;
      write_enable_data_log_force[2775] <= 1'h0;
      write_enable_data_log_force[2776] <= 1'h0;
      write_enable_data_log_force[2777] <= 1'h0;
      write_enable_data_log_force[2778] <= 1'h0;
      write_enable_data_log_force[2779] <= 1'h0;
      write_enable_data_log_force[2780] <= 1'h0;
      write_enable_data_log_force[2781] <= 1'h0;
      write_enable_data_log_force[2782] <= 1'h0;
      write_enable_data_log_force[2783] <= 1'h0;
      write_enable_data_log_force[2784] <= 1'h0;
      write_enable_data_log_force[2785] <= 1'h0;
      write_enable_data_log_force[2786] <= 1'h0;
      write_enable_data_log_force[2787] <= 1'h0;
      write_enable_data_log_force[2788] <= 1'h0;
      write_enable_data_log_force[2789] <= 1'h0;
      write_enable_data_log_force[2790] <= 1'h0;
      write_enable_data_log_force[2791] <= 1'h0;
      write_enable_data_log_force[2792] <= 1'h0;
      write_enable_data_log_force[2793] <= 1'h0;
      write_enable_data_log_force[2794] <= 1'h0;
      write_enable_data_log_force[2795] <= 1'h0;
      write_enable_data_log_force[2796] <= 1'h0;
      write_enable_data_log_force[2797] <= 1'h0;
      write_enable_data_log_force[2798] <= 1'h0;
      write_enable_data_log_force[2799] <= 1'h0;
      write_enable_data_log_force[2800] <= 1'h0;
      write_enable_data_log_force[2801] <= 1'h0;
      write_enable_data_log_force[2802] <= 1'h0;
      write_enable_data_log_force[2803] <= 1'h0;
      write_enable_data_log_force[2804] <= 1'h0;
      write_enable_data_log_force[2805] <= 1'h0;
      write_enable_data_log_force[2806] <= 1'h0;
      write_enable_data_log_force[2807] <= 1'h0;
      write_enable_data_log_force[2808] <= 1'h0;
      write_enable_data_log_force[2809] <= 1'h0;
      write_enable_data_log_force[2810] <= 1'h0;
      write_enable_data_log_force[2811] <= 1'h0;
      write_enable_data_log_force[2812] <= 1'h0;
      write_enable_data_log_force[2813] <= 1'h0;
      write_enable_data_log_force[2814] <= 1'h0;
      write_enable_data_log_force[2815] <= 1'h0;
      write_enable_data_log_force[2816] <= 1'h0;
      write_enable_data_log_force[2817] <= 1'h0;
      write_enable_data_log_force[2818] <= 1'h0;
      write_enable_data_log_force[2819] <= 1'h0;
      write_enable_data_log_force[2820] <= 1'h0;
      write_enable_data_log_force[2821] <= 1'h0;
      write_enable_data_log_force[2822] <= 1'h0;
      write_enable_data_log_force[2823] <= 1'h0;
      write_enable_data_log_force[2824] <= 1'h0;
      write_enable_data_log_force[2825] <= 1'h0;
      write_enable_data_log_force[2826] <= 1'h0;
      write_enable_data_log_force[2827] <= 1'h0;
      write_enable_data_log_force[2828] <= 1'h0;
      write_enable_data_log_force[2829] <= 1'h0;
      write_enable_data_log_force[2830] <= 1'h0;
      write_enable_data_log_force[2831] <= 1'h0;
      write_enable_data_log_force[2832] <= 1'h0;
      write_enable_data_log_force[2833] <= 1'h0;
      write_enable_data_log_force[2834] <= 1'h0;
      write_enable_data_log_force[2835] <= 1'h0;
      write_enable_data_log_force[2836] <= 1'h0;
      write_enable_data_log_force[2837] <= 1'h0;
      write_enable_data_log_force[2838] <= 1'h0;
      write_enable_data_log_force[2839] <= 1'h0;
      write_enable_data_log_force[2840] <= 1'h0;
      write_enable_data_log_force[2841] <= 1'h0;
      write_enable_data_log_force[2842] <= 1'h0;
      write_enable_data_log_force[2843] <= 1'h0;
      write_enable_data_log_force[2844] <= 1'h0;
      write_enable_data_log_force[2845] <= 1'h0;
      write_enable_data_log_force[2846] <= 1'h0;
      write_enable_data_log_force[2847] <= 1'h0;
      write_enable_data_log_force[2848] <= 1'h0;
      write_enable_data_log_force[2849] <= 1'h0;
      write_enable_data_log_force[2850] <= 1'h0;
      write_enable_data_log_force[2851] <= 1'h0;
      write_enable_data_log_force[2852] <= 1'h0;
      write_enable_data_log_force[2853] <= 1'h0;
      write_enable_data_log_force[2854] <= 1'h0;
      write_enable_data_log_force[2855] <= 1'h0;
      write_enable_data_log_force[2856] <= 1'h0;
      write_enable_data_log_force[2857] <= 1'h0;
      write_enable_data_log_force[2858] <= 1'h0;
      write_enable_data_log_force[2859] <= 1'h0;
      write_enable_data_log_force[2860] <= 1'h0;
      write_enable_data_log_force[2861] <= 1'h0;
      write_enable_data_log_force[2862] <= 1'h0;
      write_enable_data_log_force[2863] <= 1'h0;
      write_enable_data_log_force[2864] <= 1'h0;
      write_enable_data_log_force[2865] <= 1'h0;
      write_enable_data_log_force[2866] <= 1'h0;
      write_enable_data_log_force[2867] <= 1'h0;
      write_enable_data_log_force[2868] <= 1'h0;
      write_enable_data_log_force[2869] <= 1'h0;
      write_enable_data_log_force[2870] <= 1'h0;
      write_enable_data_log_force[2871] <= 1'h0;
      write_enable_data_log_force[2872] <= 1'h0;
      write_enable_data_log_force[2873] <= 1'h0;
      write_enable_data_log_force[2874] <= 1'h0;
      write_enable_data_log_force[2875] <= 1'h0;
      write_enable_data_log_force[2876] <= 1'h0;
      write_enable_data_log_force[2877] <= 1'h0;
      write_enable_data_log_force[2878] <= 1'h0;
      write_enable_data_log_force[2879] <= 1'h0;
      write_enable_data_log_force[2880] <= 1'h0;
      write_enable_data_log_force[2881] <= 1'h0;
      write_enable_data_log_force[2882] <= 1'h0;
      write_enable_data_log_force[2883] <= 1'h0;
      write_enable_data_log_force[2884] <= 1'h0;
      write_enable_data_log_force[2885] <= 1'h0;
      write_enable_data_log_force[2886] <= 1'h0;
      write_enable_data_log_force[2887] <= 1'h0;
      write_enable_data_log_force[2888] <= 1'h0;
      write_enable_data_log_force[2889] <= 1'h0;
      write_enable_data_log_force[2890] <= 1'h0;
      write_enable_data_log_force[2891] <= 1'h0;
      write_enable_data_log_force[2892] <= 1'h0;
      write_enable_data_log_force[2893] <= 1'h0;
      write_enable_data_log_force[2894] <= 1'h0;
      write_enable_data_log_force[2895] <= 1'h0;
      write_enable_data_log_force[2896] <= 1'h0;
      write_enable_data_log_force[2897] <= 1'h0;
      write_enable_data_log_force[2898] <= 1'h0;
      write_enable_data_log_force[2899] <= 1'h0;
      write_enable_data_log_force[2900] <= 1'h0;
      write_enable_data_log_force[2901] <= 1'h0;
      write_enable_data_log_force[2902] <= 1'h0;
      write_enable_data_log_force[2903] <= 1'h0;
      write_enable_data_log_force[2904] <= 1'h0;
      write_enable_data_log_force[2905] <= 1'h0;
      write_enable_data_log_force[2906] <= 1'h0;
      write_enable_data_log_force[2907] <= 1'h0;
      write_enable_data_log_force[2908] <= 1'h0;
      write_enable_data_log_force[2909] <= 1'h0;
      write_enable_data_log_force[2910] <= 1'h0;
      write_enable_data_log_force[2911] <= 1'h0;
      write_enable_data_log_force[2912] <= 1'h0;
      write_enable_data_log_force[2913] <= 1'h0;
      write_enable_data_log_force[2914] <= 1'h0;
      write_enable_data_log_force[2915] <= 1'h0;
      write_enable_data_log_force[2916] <= 1'h0;
      write_enable_data_log_force[2917] <= 1'h0;
      write_enable_data_log_force[2918] <= 1'h0;
      write_enable_data_log_force[2919] <= 1'h0;
      write_enable_data_log_force[2920] <= 1'h0;
      write_enable_data_log_force[2921] <= 1'h0;
      write_enable_data_log_force[2922] <= 1'h0;
      write_enable_data_log_force[2923] <= 1'h0;
      write_enable_data_log_force[2924] <= 1'h0;
      write_enable_data_log_force[2925] <= 1'h0;
      write_enable_data_log_force[2926] <= 1'h0;
      write_enable_data_log_force[2927] <= 1'h0;
      write_enable_data_log_force[2928] <= 1'h0;
      write_enable_data_log_force[2929] <= 1'h0;
      write_enable_data_log_force[2930] <= 1'h0;
      write_enable_data_log_force[2931] <= 1'h0;
      write_enable_data_log_force[2932] <= 1'h0;
      write_enable_data_log_force[2933] <= 1'h0;
      write_enable_data_log_force[2934] <= 1'h0;
      write_enable_data_log_force[2935] <= 1'h0;
      write_enable_data_log_force[2936] <= 1'h0;
      write_enable_data_log_force[2937] <= 1'h0;
      write_enable_data_log_force[2938] <= 1'h0;
      write_enable_data_log_force[2939] <= 1'h0;
      write_enable_data_log_force[2940] <= 1'h0;
      write_enable_data_log_force[2941] <= 1'h0;
      write_enable_data_log_force[2942] <= 1'h0;
      write_enable_data_log_force[2943] <= 1'h0;
      write_enable_data_log_force[2944] <= 1'h0;
      write_enable_data_log_force[2945] <= 1'h0;
      write_enable_data_log_force[2946] <= 1'h0;
      write_enable_data_log_force[2947] <= 1'h0;
      write_enable_data_log_force[2948] <= 1'h0;
      write_enable_data_log_force[2949] <= 1'h0;
      write_enable_data_log_force[2950] <= 1'h0;
      write_enable_data_log_force[2951] <= 1'h0;
      write_enable_data_log_force[2952] <= 1'h0;
      write_enable_data_log_force[2953] <= 1'h0;
      write_enable_data_log_force[2954] <= 1'h0;
      write_enable_data_log_force[2955] <= 1'h0;
      write_enable_data_log_force[2956] <= 1'h0;
      write_enable_data_log_force[2957] <= 1'h0;
      write_enable_data_log_force[2958] <= 1'h0;
      write_enable_data_log_force[2959] <= 1'h0;
      write_enable_data_log_force[2960] <= 1'h0;
      write_enable_data_log_force[2961] <= 1'h0;
      write_enable_data_log_force[2962] <= 1'h0;
      write_enable_data_log_force[2963] <= 1'h0;
      write_enable_data_log_force[2964] <= 1'h0;
      write_enable_data_log_force[2965] <= 1'h0;
      write_enable_data_log_force[2966] <= 1'h0;
      write_enable_data_log_force[2967] <= 1'h0;
      write_enable_data_log_force[2968] <= 1'h0;
      write_enable_data_log_force[2969] <= 1'h0;
      write_enable_data_log_force[2970] <= 1'h0;
      write_enable_data_log_force[2971] <= 1'h0;
      write_enable_data_log_force[2972] <= 1'h0;
      write_enable_data_log_force[2973] <= 1'h0;
      write_enable_data_log_force[2974] <= 1'h0;
      write_enable_data_log_force[2975] <= 1'h0;
      write_enable_data_log_force[2976] <= 1'h0;
      write_enable_data_log_force[2977] <= 1'h0;
      write_enable_data_log_force[2978] <= 1'h0;
      write_enable_data_log_force[2979] <= 1'h0;
      write_enable_data_log_force[2980] <= 1'h0;
      write_enable_data_log_force[2981] <= 1'h0;
      write_enable_data_log_force[2982] <= 1'h0;
      write_enable_data_log_force[2983] <= 1'h0;
      write_enable_data_log_force[2984] <= 1'h0;
      write_enable_data_log_force[2985] <= 1'h0;
      write_enable_data_log_force[2986] <= 1'h0;
      write_enable_data_log_force[2987] <= 1'h0;
      write_enable_data_log_force[2988] <= 1'h0;
      write_enable_data_log_force[2989] <= 1'h0;
      write_enable_data_log_force[2990] <= 1'h0;
      write_enable_data_log_force[2991] <= 1'h0;
      write_enable_data_log_force[2992] <= 1'h0;
      write_enable_data_log_force[2993] <= 1'h0;
      write_enable_data_log_force[2994] <= 1'h0;
      write_enable_data_log_force[2995] <= 1'h0;
      write_enable_data_log_force[2996] <= 1'h0;
      write_enable_data_log_force[2997] <= 1'h0;
      write_enable_data_log_force[2998] <= 1'h0;
      write_enable_data_log_force[2999] <= 1'h0;
      write_enable_data_log_force[3000] <= 1'h0;
      write_enable_data_log_force[3001] <= 1'h0;
      write_enable_data_log_force[3002] <= 1'h0;
      write_enable_data_log_force[3003] <= 1'h0;
      write_enable_data_log_force[3004] <= 1'h0;
      write_enable_data_log_force[3005] <= 1'h0;
      write_enable_data_log_force[3006] <= 1'h0;
      write_enable_data_log_force[3007] <= 1'h0;
      write_enable_data_log_force[3008] <= 1'h0;
      write_enable_data_log_force[3009] <= 1'h0;
      write_enable_data_log_force[3010] <= 1'h0;
      write_enable_data_log_force[3011] <= 1'h0;
      write_enable_data_log_force[3012] <= 1'h0;
      write_enable_data_log_force[3013] <= 1'h0;
      write_enable_data_log_force[3014] <= 1'h0;
      write_enable_data_log_force[3015] <= 1'h0;
      write_enable_data_log_force[3016] <= 1'h0;
      write_enable_data_log_force[3017] <= 1'h0;
      write_enable_data_log_force[3018] <= 1'h0;
      write_enable_data_log_force[3019] <= 1'h0;
      write_enable_data_log_force[3020] <= 1'h0;
      write_enable_data_log_force[3021] <= 1'h0;
      write_enable_data_log_force[3022] <= 1'h0;
      write_enable_data_log_force[3023] <= 1'h0;
      write_enable_data_log_force[3024] <= 1'h0;
      write_enable_data_log_force[3025] <= 1'h0;
      write_enable_data_log_force[3026] <= 1'h0;
      write_enable_data_log_force[3027] <= 1'h0;
      write_enable_data_log_force[3028] <= 1'h0;
      write_enable_data_log_force[3029] <= 1'h0;
      write_enable_data_log_force[3030] <= 1'h0;
      write_enable_data_log_force[3031] <= 1'h0;
      write_enable_data_log_force[3032] <= 1'h0;
      write_enable_data_log_force[3033] <= 1'h0;
      write_enable_data_log_force[3034] <= 1'h0;
      write_enable_data_log_force[3035] <= 1'h0;
      write_enable_data_log_force[3036] <= 1'h0;
      write_enable_data_log_force[3037] <= 1'h0;
      write_enable_data_log_force[3038] <= 1'h0;
      write_enable_data_log_force[3039] <= 1'h0;
      write_enable_data_log_force[3040] <= 1'h0;
      write_enable_data_log_force[3041] <= 1'h0;
      write_enable_data_log_force[3042] <= 1'h0;
      write_enable_data_log_force[3043] <= 1'h0;
      write_enable_data_log_force[3044] <= 1'h0;
      write_enable_data_log_force[3045] <= 1'h0;
      write_enable_data_log_force[3046] <= 1'h0;
      write_enable_data_log_force[3047] <= 1'h0;
      write_enable_data_log_force[3048] <= 1'h0;
      write_enable_data_log_force[3049] <= 1'h0;
      write_enable_data_log_force[3050] <= 1'h0;
      write_enable_data_log_force[3051] <= 1'h0;
      write_enable_data_log_force[3052] <= 1'h0;
      write_enable_data_log_force[3053] <= 1'h0;
      write_enable_data_log_force[3054] <= 1'h0;
      write_enable_data_log_force[3055] <= 1'h0;
      write_enable_data_log_force[3056] <= 1'h0;
      write_enable_data_log_force[3057] <= 1'h0;
      write_enable_data_log_force[3058] <= 1'h0;
      write_enable_data_log_force[3059] <= 1'h0;
      write_enable_data_log_force[3060] <= 1'h0;
      write_enable_data_log_force[3061] <= 1'h0;
      write_enable_data_log_force[3062] <= 1'h0;
      write_enable_data_log_force[3063] <= 1'h0;
      write_enable_data_log_force[3064] <= 1'h0;
      write_enable_data_log_force[3065] <= 1'h0;
      write_enable_data_log_force[3066] <= 1'h0;
      write_enable_data_log_force[3067] <= 1'h0;
      write_enable_data_log_force[3068] <= 1'h0;
      write_enable_data_log_force[3069] <= 1'h0;
      write_enable_data_log_force[3070] <= 1'h0;
      write_enable_data_log_force[3071] <= 1'h0;
      write_enable_data_log_force[3072] <= 1'h0;
      write_enable_data_log_force[3073] <= 1'h0;
      write_enable_data_log_force[3074] <= 1'h0;
      write_enable_data_log_force[3075] <= 1'h0;
      write_enable_data_log_force[3076] <= 1'h0;
      write_enable_data_log_force[3077] <= 1'h0;
      write_enable_data_log_force[3078] <= 1'h0;
      write_enable_data_log_force[3079] <= 1'h0;
      write_enable_data_log_force[3080] <= 1'h0;
      write_enable_data_log_force[3081] <= 1'h0;
      write_enable_data_log_force[3082] <= 1'h0;
      write_enable_data_log_force[3083] <= 1'h0;
      write_enable_data_log_force[3084] <= 1'h0;
      write_enable_data_log_force[3085] <= 1'h0;
      write_enable_data_log_force[3086] <= 1'h0;
      write_enable_data_log_force[3087] <= 1'h0;
      write_enable_data_log_force[3088] <= 1'h0;
      write_enable_data_log_force[3089] <= 1'h0;
      write_enable_data_log_force[3090] <= 1'h0;
      write_enable_data_log_force[3091] <= 1'h0;
      write_enable_data_log_force[3092] <= 1'h0;
      write_enable_data_log_force[3093] <= 1'h0;
      write_enable_data_log_force[3094] <= 1'h0;
      write_enable_data_log_force[3095] <= 1'h0;
      write_enable_data_log_force[3096] <= 1'h0;
      write_enable_data_log_force[3097] <= 1'h0;
      write_enable_data_log_force[3098] <= 1'h0;
      write_enable_data_log_force[3099] <= 1'h0;
      write_enable_data_log_force[3100] <= 1'h0;
      write_enable_data_log_force[3101] <= 1'h0;
      write_enable_data_log_force[3102] <= 1'h0;
      write_enable_data_log_force[3103] <= 1'h0;
      write_enable_data_log_force[3104] <= 1'h0;
      write_enable_data_log_force[3105] <= 1'h0;
      write_enable_data_log_force[3106] <= 1'h0;
      write_enable_data_log_force[3107] <= 1'h0;
      write_enable_data_log_force[3108] <= 1'h0;
      write_enable_data_log_force[3109] <= 1'h0;
      write_enable_data_log_force[3110] <= 1'h0;
      write_enable_data_log_force[3111] <= 1'h0;
      write_enable_data_log_force[3112] <= 1'h0;
      write_enable_data_log_force[3113] <= 1'h0;
      write_enable_data_log_force[3114] <= 1'h0;
      write_enable_data_log_force[3115] <= 1'h0;
      write_enable_data_log_force[3116] <= 1'h0;
      write_enable_data_log_force[3117] <= 1'h0;
      write_enable_data_log_force[3118] <= 1'h0;
      write_enable_data_log_force[3119] <= 1'h0;
      write_enable_data_log_force[3120] <= 1'h0;
      write_enable_data_log_force[3121] <= 1'h0;
      write_enable_data_log_force[3122] <= 1'h0;
      write_enable_data_log_force[3123] <= 1'h0;
      write_enable_data_log_force[3124] <= 1'h0;
      write_enable_data_log_force[3125] <= 1'h0;
      write_enable_data_log_force[3126] <= 1'h0;
      write_enable_data_log_force[3127] <= 1'h0;
      write_enable_data_log_force[3128] <= 1'h0;
      write_enable_data_log_force[3129] <= 1'h0;
      write_enable_data_log_force[3130] <= 1'h0;
      write_enable_data_log_force[3131] <= 1'h0;
      write_enable_data_log_force[3132] <= 1'h0;
      write_enable_data_log_force[3133] <= 1'h0;
      write_enable_data_log_force[3134] <= 1'h0;
      write_enable_data_log_force[3135] <= 1'h0;
      write_enable_data_log_force[3136] <= 1'h0;
      write_enable_data_log_force[3137] <= 1'h0;
      write_enable_data_log_force[3138] <= 1'h0;
      write_enable_data_log_force[3139] <= 1'h0;
      write_enable_data_log_force[3140] <= 1'h0;
      write_enable_data_log_force[3141] <= 1'h0;
      write_enable_data_log_force[3142] <= 1'h0;
      write_enable_data_log_force[3143] <= 1'h0;
      write_enable_data_log_force[3144] <= 1'h0;
      write_enable_data_log_force[3145] <= 1'h0;
      write_enable_data_log_force[3146] <= 1'h0;
      write_enable_data_log_force[3147] <= 1'h0;
      write_enable_data_log_force[3148] <= 1'h0;
      write_enable_data_log_force[3149] <= 1'h0;
      write_enable_data_log_force[3150] <= 1'h0;
      write_enable_data_log_force[3151] <= 1'h0;
      write_enable_data_log_force[3152] <= 1'h0;
      write_enable_data_log_force[3153] <= 1'h0;
      write_enable_data_log_force[3154] <= 1'h0;
      write_enable_data_log_force[3155] <= 1'h0;
      write_enable_data_log_force[3156] <= 1'h0;
      write_enable_data_log_force[3157] <= 1'h0;
      write_enable_data_log_force[3158] <= 1'h0;
      write_enable_data_log_force[3159] <= 1'h0;
      write_enable_data_log_force[3160] <= 1'h0;
      write_enable_data_log_force[3161] <= 1'h0;
      write_enable_data_log_force[3162] <= 1'h0;
      write_enable_data_log_force[3163] <= 1'h0;
      write_enable_data_log_force[3164] <= 1'h0;
      write_enable_data_log_force[3165] <= 1'h0;
      write_enable_data_log_force[3166] <= 1'h0;
      write_enable_data_log_force[3167] <= 1'h0;
      write_enable_data_log_force[3168] <= 1'h0;
      write_enable_data_log_force[3169] <= 1'h0;
      write_enable_data_log_force[3170] <= 1'h0;
      write_enable_data_log_force[3171] <= 1'h0;
      write_enable_data_log_force[3172] <= 1'h0;
      write_enable_data_log_force[3173] <= 1'h0;
      write_enable_data_log_force[3174] <= 1'h0;
      write_enable_data_log_force[3175] <= 1'h0;
      write_enable_data_log_force[3176] <= 1'h0;
      write_enable_data_log_force[3177] <= 1'h0;
      write_enable_data_log_force[3178] <= 1'h0;
      write_enable_data_log_force[3179] <= 1'h0;
      write_enable_data_log_force[3180] <= 1'h0;
      write_enable_data_log_force[3181] <= 1'h0;
      write_enable_data_log_force[3182] <= 1'h0;
      write_enable_data_log_force[3183] <= 1'h0;
      write_enable_data_log_force[3184] <= 1'h0;
      write_enable_data_log_force[3185] <= 1'h0;
      write_enable_data_log_force[3186] <= 1'h0;
      write_enable_data_log_force[3187] <= 1'h0;
      write_enable_data_log_force[3188] <= 1'h0;
      write_enable_data_log_force[3189] <= 1'h0;
      write_enable_data_log_force[3190] <= 1'h0;
      write_enable_data_log_force[3191] <= 1'h0;
      write_enable_data_log_force[3192] <= 1'h0;
      write_enable_data_log_force[3193] <= 1'h0;
      write_enable_data_log_force[3194] <= 1'h0;
      write_enable_data_log_force[3195] <= 1'h0;
      write_enable_data_log_force[3196] <= 1'h0;
      write_enable_data_log_force[3197] <= 1'h0;
      write_enable_data_log_force[3198] <= 1'h0;
      write_enable_data_log_force[3199] <= 1'h0;
      write_enable_data_log_force[3200] <= 1'h0;
      write_enable_data_log_force[3201] <= 1'h0;
      write_enable_data_log_force[3202] <= 1'h0;
      write_enable_data_log_force[3203] <= 1'h0;
      write_enable_data_log_force[3204] <= 1'h0;
      write_enable_data_log_force[3205] <= 1'h0;
      write_enable_data_log_force[3206] <= 1'h0;
      write_enable_data_log_force[3207] <= 1'h0;
      write_enable_data_log_force[3208] <= 1'h0;
      write_enable_data_log_force[3209] <= 1'h0;
      write_enable_data_log_force[3210] <= 1'h0;
      write_enable_data_log_force[3211] <= 1'h0;
      write_enable_data_log_force[3212] <= 1'h0;
      write_enable_data_log_force[3213] <= 1'h0;
      write_enable_data_log_force[3214] <= 1'h0;
      write_enable_data_log_force[3215] <= 1'h0;
      write_enable_data_log_force[3216] <= 1'h0;
      write_enable_data_log_force[3217] <= 1'h0;
      write_enable_data_log_force[3218] <= 1'h0;
      write_enable_data_log_force[3219] <= 1'h0;
      write_enable_data_log_force[3220] <= 1'h0;
      write_enable_data_log_force[3221] <= 1'h0;
      write_enable_data_log_force[3222] <= 1'h0;
      write_enable_data_log_force[3223] <= 1'h0;
      write_enable_data_log_force[3224] <= 1'h0;
      write_enable_data_log_force[3225] <= 1'h0;
      write_enable_data_log_force[3226] <= 1'h0;
      write_enable_data_log_force[3227] <= 1'h0;
      write_enable_data_log_force[3228] <= 1'h0;
      write_enable_data_log_force[3229] <= 1'h0;
      write_enable_data_log_force[3230] <= 1'h0;
      write_enable_data_log_force[3231] <= 1'h0;
      write_enable_data_log_force[3232] <= 1'h0;
      write_enable_data_log_force[3233] <= 1'h0;
      write_enable_data_log_force[3234] <= 1'h0;
      write_enable_data_log_force[3235] <= 1'h0;
      write_enable_data_log_force[3236] <= 1'h0;
      write_enable_data_log_force[3237] <= 1'h0;
      write_enable_data_log_force[3238] <= 1'h0;
      write_enable_data_log_force[3239] <= 1'h0;
      write_enable_data_log_force[3240] <= 1'h0;
      write_enable_data_log_force[3241] <= 1'h0;
      write_enable_data_log_force[3242] <= 1'h0;
      write_enable_data_log_force[3243] <= 1'h0;
      write_enable_data_log_force[3244] <= 1'h0;
      write_enable_data_log_force[3245] <= 1'h0;
      write_enable_data_log_force[3246] <= 1'h0;
      write_enable_data_log_force[3247] <= 1'h0;
      write_enable_data_log_force[3248] <= 1'h0;
      write_enable_data_log_force[3249] <= 1'h0;
      write_enable_data_log_force[3250] <= 1'h0;
      write_enable_data_log_force[3251] <= 1'h0;
      write_enable_data_log_force[3252] <= 1'h0;
      write_enable_data_log_force[3253] <= 1'h0;
      write_enable_data_log_force[3254] <= 1'h0;
      write_enable_data_log_force[3255] <= 1'h0;
      write_enable_data_log_force[3256] <= 1'h0;
      write_enable_data_log_force[3257] <= 1'h0;
      write_enable_data_log_force[3258] <= 1'h0;
      write_enable_data_log_force[3259] <= 1'h0;
      write_enable_data_log_force[3260] <= 1'h0;
      write_enable_data_log_force[3261] <= 1'h0;
      write_enable_data_log_force[3262] <= 1'h0;
      write_enable_data_log_force[3263] <= 1'h0;
      write_enable_data_log_force[3264] <= 1'h0;
      write_enable_data_log_force[3265] <= 1'h0;
      write_enable_data_log_force[3266] <= 1'h0;
      write_enable_data_log_force[3267] <= 1'h0;
      write_enable_data_log_force[3268] <= 1'h0;
      write_enable_data_log_force[3269] <= 1'h0;
      write_enable_data_log_force[3270] <= 1'h0;
      write_enable_data_log_force[3271] <= 1'h0;
      write_enable_data_log_force[3272] <= 1'h0;
      write_enable_data_log_force[3273] <= 1'h0;
      write_enable_data_log_force[3274] <= 1'h0;
      write_enable_data_log_force[3275] <= 1'h0;
      write_enable_data_log_force[3276] <= 1'h0;
      write_enable_data_log_force[3277] <= 1'h0;
      write_enable_data_log_force[3278] <= 1'h0;
      write_enable_data_log_force[3279] <= 1'h0;
      write_enable_data_log_force[3280] <= 1'h0;
      write_enable_data_log_force[3281] <= 1'h0;
      write_enable_data_log_force[3282] <= 1'h0;
      write_enable_data_log_force[3283] <= 1'h0;
      write_enable_data_log_force[3284] <= 1'h0;
      write_enable_data_log_force[3285] <= 1'h0;
      write_enable_data_log_force[3286] <= 1'h0;
      write_enable_data_log_force[3287] <= 1'h0;
      write_enable_data_log_force[3288] <= 1'h0;
      write_enable_data_log_force[3289] <= 1'h0;
      write_enable_data_log_force[3290] <= 1'h0;
      write_enable_data_log_force[3291] <= 1'h0;
      write_enable_data_log_force[3292] <= 1'h0;
      write_enable_data_log_force[3293] <= 1'h0;
      write_enable_data_log_force[3294] <= 1'h0;
      write_enable_data_log_force[3295] <= 1'h0;
      write_enable_data_log_force[3296] <= 1'h0;
      write_enable_data_log_force[3297] <= 1'h0;
      write_enable_data_log_force[3298] <= 1'h0;
      write_enable_data_log_force[3299] <= 1'h0;
      write_enable_data_log_force[3300] <= 1'h0;
      write_enable_data_log_force[3301] <= 1'h0;
      write_enable_data_log_force[3302] <= 1'h0;
      write_enable_data_log_force[3303] <= 1'h0;
      write_enable_data_log_force[3304] <= 1'h0;
      write_enable_data_log_force[3305] <= 1'h0;
      write_enable_data_log_force[3306] <= 1'h0;
      write_enable_data_log_force[3307] <= 1'h0;
      write_enable_data_log_force[3308] <= 1'h0;
      write_enable_data_log_force[3309] <= 1'h0;
      write_enable_data_log_force[3310] <= 1'h0;
      write_enable_data_log_force[3311] <= 1'h0;
      write_enable_data_log_force[3312] <= 1'h0;
      write_enable_data_log_force[3313] <= 1'h0;
      write_enable_data_log_force[3314] <= 1'h0;
      write_enable_data_log_force[3315] <= 1'h0;
      write_enable_data_log_force[3316] <= 1'h0;
      write_enable_data_log_force[3317] <= 1'h0;
      write_enable_data_log_force[3318] <= 1'h0;
      write_enable_data_log_force[3319] <= 1'h0;
      write_enable_data_log_force[3320] <= 1'h0;
      write_enable_data_log_force[3321] <= 1'h0;
      write_enable_data_log_force[3322] <= 1'h0;
      write_enable_data_log_force[3323] <= 1'h0;
      write_enable_data_log_force[3324] <= 1'h0;
      write_enable_data_log_force[3325] <= 1'h0;
      write_enable_data_log_force[3326] <= 1'h0;
      write_enable_data_log_force[3327] <= 1'h0;
      write_enable_data_log_force[3328] <= 1'h0;
      write_enable_data_log_force[3329] <= 1'h0;
      write_enable_data_log_force[3330] <= 1'h0;
      write_enable_data_log_force[3331] <= 1'h0;
      write_enable_data_log_force[3332] <= 1'h0;
      write_enable_data_log_force[3333] <= 1'h0;
      write_enable_data_log_force[3334] <= 1'h0;
      write_enable_data_log_force[3335] <= 1'h0;
      write_enable_data_log_force[3336] <= 1'h0;
      write_enable_data_log_force[3337] <= 1'h0;
      write_enable_data_log_force[3338] <= 1'h0;
      write_enable_data_log_force[3339] <= 1'h0;
      write_enable_data_log_force[3340] <= 1'h0;
      write_enable_data_log_force[3341] <= 1'h0;
      write_enable_data_log_force[3342] <= 1'h0;
      write_enable_data_log_force[3343] <= 1'h0;
      write_enable_data_log_force[3344] <= 1'h0;
      write_enable_data_log_force[3345] <= 1'h0;
      write_enable_data_log_force[3346] <= 1'h0;
      write_enable_data_log_force[3347] <= 1'h0;
      write_enable_data_log_force[3348] <= 1'h0;
      write_enable_data_log_force[3349] <= 1'h0;
      write_enable_data_log_force[3350] <= 1'h0;
      write_enable_data_log_force[3351] <= 1'h0;
      write_enable_data_log_force[3352] <= 1'h0;
      write_enable_data_log_force[3353] <= 1'h0;
      write_enable_data_log_force[3354] <= 1'h0;
      write_enable_data_log_force[3355] <= 1'h0;
      write_enable_data_log_force[3356] <= 1'h0;
      write_enable_data_log_force[3357] <= 1'h0;
      write_enable_data_log_force[3358] <= 1'h0;
      write_enable_data_log_force[3359] <= 1'h0;
      write_enable_data_log_force[3360] <= 1'h0;
      write_enable_data_log_force[3361] <= 1'h0;
      write_enable_data_log_force[3362] <= 1'h0;
      write_enable_data_log_force[3363] <= 1'h0;
      write_enable_data_log_force[3364] <= 1'h0;
      write_enable_data_log_force[3365] <= 1'h0;
      write_enable_data_log_force[3366] <= 1'h0;
      write_enable_data_log_force[3367] <= 1'h0;
      write_enable_data_log_force[3368] <= 1'h0;
      write_enable_data_log_force[3369] <= 1'h0;
      write_enable_data_log_force[3370] <= 1'h0;
      write_enable_data_log_force[3371] <= 1'h0;
      write_enable_data_log_force[3372] <= 1'h0;
      write_enable_data_log_force[3373] <= 1'h0;
      write_enable_data_log_force[3374] <= 1'h0;
      write_enable_data_log_force[3375] <= 1'h0;
      write_enable_data_log_force[3376] <= 1'h0;
      write_enable_data_log_force[3377] <= 1'h0;
      write_enable_data_log_force[3378] <= 1'h0;
      write_enable_data_log_force[3379] <= 1'h0;
      write_enable_data_log_force[3380] <= 1'h0;
      write_enable_data_log_force[3381] <= 1'h0;
      write_enable_data_log_force[3382] <= 1'h0;
      write_enable_data_log_force[3383] <= 1'h0;
      write_enable_data_log_force[3384] <= 1'h0;
      write_enable_data_log_force[3385] <= 1'h0;
      write_enable_data_log_force[3386] <= 1'h0;
      write_enable_data_log_force[3387] <= 1'h0;
      write_enable_data_log_force[3388] <= 1'h0;
      write_enable_data_log_force[3389] <= 1'h0;
      write_enable_data_log_force[3390] <= 1'h0;
      write_enable_data_log_force[3391] <= 1'h0;
      write_enable_data_log_force[3392] <= 1'h0;
      write_enable_data_log_force[3393] <= 1'h0;
      write_enable_data_log_force[3394] <= 1'h0;
      write_enable_data_log_force[3395] <= 1'h0;
      write_enable_data_log_force[3396] <= 1'h0;
      write_enable_data_log_force[3397] <= 1'h0;
      write_enable_data_log_force[3398] <= 1'h0;
      write_enable_data_log_force[3399] <= 1'h0;
      write_enable_data_log_force[3400] <= 1'h0;
      write_enable_data_log_force[3401] <= 1'h0;
      write_enable_data_log_force[3402] <= 1'h0;
      write_enable_data_log_force[3403] <= 1'h0;
      write_enable_data_log_force[3404] <= 1'h0;
      write_enable_data_log_force[3405] <= 1'h0;
      write_enable_data_log_force[3406] <= 1'h0;
      write_enable_data_log_force[3407] <= 1'h0;
      write_enable_data_log_force[3408] <= 1'h0;
      write_enable_data_log_force[3409] <= 1'h0;
      write_enable_data_log_force[3410] <= 1'h0;
      write_enable_data_log_force[3411] <= 1'h0;
      write_enable_data_log_force[3412] <= 1'h0;
      write_enable_data_log_force[3413] <= 1'h0;
      write_enable_data_log_force[3414] <= 1'h0;
      write_enable_data_log_force[3415] <= 1'h0;
      write_enable_data_log_force[3416] <= 1'h0;
      write_enable_data_log_force[3417] <= 1'h0;
      write_enable_data_log_force[3418] <= 1'h0;
      write_enable_data_log_force[3419] <= 1'h0;
      write_enable_data_log_force[3420] <= 1'h0;
      write_enable_data_log_force[3421] <= 1'h0;
      write_enable_data_log_force[3422] <= 1'h0;
      write_enable_data_log_force[3423] <= 1'h0;
      write_enable_data_log_force[3424] <= 1'h0;
      write_enable_data_log_force[3425] <= 1'h0;
      write_enable_data_log_force[3426] <= 1'h0;
      write_enable_data_log_force[3427] <= 1'h0;
      write_enable_data_log_force[3428] <= 1'h0;
      write_enable_data_log_force[3429] <= 1'h0;
      write_enable_data_log_force[3430] <= 1'h0;
      write_enable_data_log_force[3431] <= 1'h0;
      write_enable_data_log_force[3432] <= 1'h0;
      write_enable_data_log_force[3433] <= 1'h0;
      write_enable_data_log_force[3434] <= 1'h0;
      write_enable_data_log_force[3435] <= 1'h0;
      write_enable_data_log_force[3436] <= 1'h0;
      write_enable_data_log_force[3437] <= 1'h0;
      write_enable_data_log_force[3438] <= 1'h0;
      write_enable_data_log_force[3439] <= 1'h0;
      write_enable_data_log_force[3440] <= 1'h0;
      write_enable_data_log_force[3441] <= 1'h0;
      write_enable_data_log_force[3442] <= 1'h0;
      write_enable_data_log_force[3443] <= 1'h0;
      write_enable_data_log_force[3444] <= 1'h0;
      write_enable_data_log_force[3445] <= 1'h0;
      write_enable_data_log_force[3446] <= 1'h0;
      write_enable_data_log_force[3447] <= 1'h0;
      write_enable_data_log_force[3448] <= 1'h0;
      write_enable_data_log_force[3449] <= 1'h0;
      write_enable_data_log_force[3450] <= 1'h0;
      write_enable_data_log_force[3451] <= 1'h0;
      write_enable_data_log_force[3452] <= 1'h0;
      write_enable_data_log_force[3453] <= 1'h0;
      write_enable_data_log_force[3454] <= 1'h0;
      write_enable_data_log_force[3455] <= 1'h0;
      write_enable_data_log_force[3456] <= 1'h0;
      write_enable_data_log_force[3457] <= 1'h0;
      write_enable_data_log_force[3458] <= 1'h0;
      write_enable_data_log_force[3459] <= 1'h0;
      write_enable_data_log_force[3460] <= 1'h0;
      write_enable_data_log_force[3461] <= 1'h0;
      write_enable_data_log_force[3462] <= 1'h0;
      write_enable_data_log_force[3463] <= 1'h0;
      write_enable_data_log_force[3464] <= 1'h0;
      write_enable_data_log_force[3465] <= 1'h0;
      write_enable_data_log_force[3466] <= 1'h0;
      write_enable_data_log_force[3467] <= 1'h0;
      write_enable_data_log_force[3468] <= 1'h0;
      write_enable_data_log_force[3469] <= 1'h0;
      write_enable_data_log_force[3470] <= 1'h0;
      write_enable_data_log_force[3471] <= 1'h0;
      write_enable_data_log_force[3472] <= 1'h0;
      write_enable_data_log_force[3473] <= 1'h0;
      write_enable_data_log_force[3474] <= 1'h0;
      write_enable_data_log_force[3475] <= 1'h0;
      write_enable_data_log_force[3476] <= 1'h0;
      write_enable_data_log_force[3477] <= 1'h0;
      write_enable_data_log_force[3478] <= 1'h0;
      write_enable_data_log_force[3479] <= 1'h0;
      write_enable_data_log_force[3480] <= 1'h0;
      write_enable_data_log_force[3481] <= 1'h0;
      write_enable_data_log_force[3482] <= 1'h0;
      write_enable_data_log_force[3483] <= 1'h0;
      write_enable_data_log_force[3484] <= 1'h0;
      write_enable_data_log_force[3485] <= 1'h0;
      write_enable_data_log_force[3486] <= 1'h0;
      write_enable_data_log_force[3487] <= 1'h0;
      write_enable_data_log_force[3488] <= 1'h0;
      write_enable_data_log_force[3489] <= 1'h0;
      write_enable_data_log_force[3490] <= 1'h0;
      write_enable_data_log_force[3491] <= 1'h0;
      write_enable_data_log_force[3492] <= 1'h0;
      write_enable_data_log_force[3493] <= 1'h0;
      write_enable_data_log_force[3494] <= 1'h0;
      write_enable_data_log_force[3495] <= 1'h0;
      write_enable_data_log_force[3496] <= 1'h0;
      write_enable_data_log_force[3497] <= 1'h0;
      write_enable_data_log_force[3498] <= 1'h0;
      write_enable_data_log_force[3499] <= 1'h0;
      write_enable_data_log_force[3500] <= 1'h0;
      write_enable_data_log_force[3501] <= 1'h0;
      write_enable_data_log_force[3502] <= 1'h0;
      write_enable_data_log_force[3503] <= 1'h0;
      write_enable_data_log_force[3504] <= 1'h0;
      write_enable_data_log_force[3505] <= 1'h0;
      write_enable_data_log_force[3506] <= 1'h0;
      write_enable_data_log_force[3507] <= 1'h0;
      write_enable_data_log_force[3508] <= 1'h0;
      write_enable_data_log_force[3509] <= 1'h0;
      write_enable_data_log_force[3510] <= 1'h0;
      write_enable_data_log_force[3511] <= 1'h0;
      write_enable_data_log_force[3512] <= 1'h0;
      write_enable_data_log_force[3513] <= 1'h0;
      write_enable_data_log_force[3514] <= 1'h0;
      write_enable_data_log_force[3515] <= 1'h0;
      write_enable_data_log_force[3516] <= 1'h0;
      write_enable_data_log_force[3517] <= 1'h0;
      write_enable_data_log_force[3518] <= 1'h0;
      write_enable_data_log_force[3519] <= 1'h0;
      write_enable_data_log_force[3520] <= 1'h0;
      write_enable_data_log_force[3521] <= 1'h0;
      write_enable_data_log_force[3522] <= 1'h0;
      write_enable_data_log_force[3523] <= 1'h0;
      write_enable_data_log_force[3524] <= 1'h0;
      write_enable_data_log_force[3525] <= 1'h0;
      write_enable_data_log_force[3526] <= 1'h0;
      write_enable_data_log_force[3527] <= 1'h0;
      write_enable_data_log_force[3528] <= 1'h0;
      write_enable_data_log_force[3529] <= 1'h0;
      write_enable_data_log_force[3530] <= 1'h0;
      write_enable_data_log_force[3531] <= 1'h0;
      write_enable_data_log_force[3532] <= 1'h0;
      write_enable_data_log_force[3533] <= 1'h0;
      write_enable_data_log_force[3534] <= 1'h0;
      write_enable_data_log_force[3535] <= 1'h0;
      write_enable_data_log_force[3536] <= 1'h0;
      write_enable_data_log_force[3537] <= 1'h0;
      write_enable_data_log_force[3538] <= 1'h0;
      write_enable_data_log_force[3539] <= 1'h0;
      write_enable_data_log_force[3540] <= 1'h0;
      write_enable_data_log_force[3541] <= 1'h0;
      write_enable_data_log_force[3542] <= 1'h0;
      write_enable_data_log_force[3543] <= 1'h0;
      write_enable_data_log_force[3544] <= 1'h0;
      write_enable_data_log_force[3545] <= 1'h0;
      write_enable_data_log_force[3546] <= 1'h0;
      write_enable_data_log_force[3547] <= 1'h0;
      write_enable_data_log_force[3548] <= 1'h0;
      write_enable_data_log_force[3549] <= 1'h0;
      write_enable_data_log_force[3550] <= 1'h0;
      write_enable_data_log_force[3551] <= 1'h0;
      write_enable_data_log_force[3552] <= 1'h0;
      write_enable_data_log_force[3553] <= 1'h0;
      write_enable_data_log_force[3554] <= 1'h0;
      write_enable_data_log_force[3555] <= 1'h0;
      write_enable_data_log_force[3556] <= 1'h0;
      write_enable_data_log_force[3557] <= 1'h0;
      write_enable_data_log_force[3558] <= 1'h0;
      write_enable_data_log_force[3559] <= 1'h0;
      write_enable_data_log_force[3560] <= 1'h0;
      write_enable_data_log_force[3561] <= 1'h0;
      write_enable_data_log_force[3562] <= 1'h0;
      write_enable_data_log_force[3563] <= 1'h0;
      write_enable_data_log_force[3564] <= 1'h0;
      write_enable_data_log_force[3565] <= 1'h0;
      write_enable_data_log_force[3566] <= 1'h0;
      write_enable_data_log_force[3567] <= 1'h0;
      write_enable_data_log_force[3568] <= 1'h0;
      write_enable_data_log_force[3569] <= 1'h0;
      write_enable_data_log_force[3570] <= 1'h0;
      write_enable_data_log_force[3571] <= 1'h0;
      write_enable_data_log_force[3572] <= 1'h0;
      write_enable_data_log_force[3573] <= 1'h0;
      write_enable_data_log_force[3574] <= 1'h0;
      write_enable_data_log_force[3575] <= 1'h0;
      write_enable_data_log_force[3576] <= 1'h0;
      write_enable_data_log_force[3577] <= 1'h0;
      write_enable_data_log_force[3578] <= 1'h0;
      write_enable_data_log_force[3579] <= 1'h0;
      write_enable_data_log_force[3580] <= 1'h0;
      write_enable_data_log_force[3581] <= 1'h0;
      write_enable_data_log_force[3582] <= 1'h0;
      write_enable_data_log_force[3583] <= 1'h0;
      write_enable_data_log_force[3584] <= 1'h0;
      write_enable_data_log_force[3585] <= 1'h0;
      write_enable_data_log_force[3586] <= 1'h0;
      write_enable_data_log_force[3587] <= 1'h0;
      write_enable_data_log_force[3588] <= 1'h0;
      write_enable_data_log_force[3589] <= 1'h0;
      write_enable_data_log_force[3590] <= 1'h0;
      write_enable_data_log_force[3591] <= 1'h0;
      write_enable_data_log_force[3592] <= 1'h0;
      write_enable_data_log_force[3593] <= 1'h0;
      write_enable_data_log_force[3594] <= 1'h0;
      write_enable_data_log_force[3595] <= 1'h0;
      write_enable_data_log_force[3596] <= 1'h0;
      write_enable_data_log_force[3597] <= 1'h0;
      write_enable_data_log_force[3598] <= 1'h0;
      write_enable_data_log_force[3599] <= 1'h0;
      write_enable_data_log_force[3600] <= 1'h0;
      write_enable_data_log_force[3601] <= 1'h0;
      write_enable_data_log_force[3602] <= 1'h0;
      write_enable_data_log_force[3603] <= 1'h0;
      write_enable_data_log_force[3604] <= 1'h0;
      write_enable_data_log_force[3605] <= 1'h0;
      write_enable_data_log_force[3606] <= 1'h0;
      write_enable_data_log_force[3607] <= 1'h0;
      write_enable_data_log_force[3608] <= 1'h0;
      write_enable_data_log_force[3609] <= 1'h0;
      write_enable_data_log_force[3610] <= 1'h0;
      write_enable_data_log_force[3611] <= 1'h0;
      write_enable_data_log_force[3612] <= 1'h0;
      write_enable_data_log_force[3613] <= 1'h0;
      write_enable_data_log_force[3614] <= 1'h0;
      write_enable_data_log_force[3615] <= 1'h0;
      write_enable_data_log_force[3616] <= 1'h0;
      write_enable_data_log_force[3617] <= 1'h0;
      write_enable_data_log_force[3618] <= 1'h0;
      write_enable_data_log_force[3619] <= 1'h0;
      write_enable_data_log_force[3620] <= 1'h0;
      write_enable_data_log_force[3621] <= 1'h0;
      write_enable_data_log_force[3622] <= 1'h0;
      write_enable_data_log_force[3623] <= 1'h0;
      write_enable_data_log_force[3624] <= 1'h0;
      write_enable_data_log_force[3625] <= 1'h0;
      write_enable_data_log_force[3626] <= 1'h0;
      write_enable_data_log_force[3627] <= 1'h0;
      write_enable_data_log_force[3628] <= 1'h0;
      write_enable_data_log_force[3629] <= 1'h0;
      write_enable_data_log_force[3630] <= 1'h0;
      write_enable_data_log_force[3631] <= 1'h0;
      write_enable_data_log_force[3632] <= 1'h0;
      write_enable_data_log_force[3633] <= 1'h0;
      write_enable_data_log_force[3634] <= 1'h0;
      write_enable_data_log_force[3635] <= 1'h0;
      write_enable_data_log_force[3636] <= 1'h0;
      write_enable_data_log_force[3637] <= 1'h0;
      write_enable_data_log_force[3638] <= 1'h0;
      write_enable_data_log_force[3639] <= 1'h0;
      write_enable_data_log_force[3640] <= 1'h0;
      write_enable_data_log_force[3641] <= 1'h0;
      write_enable_data_log_force[3642] <= 1'h0;
      write_enable_data_log_force[3643] <= 1'h0;
      write_enable_data_log_force[3644] <= 1'h0;
      write_enable_data_log_force[3645] <= 1'h0;
      write_enable_data_log_force[3646] <= 1'h0;
      write_enable_data_log_force[3647] <= 1'h0;
      write_enable_data_log_force[3648] <= 1'h0;
      write_enable_data_log_force[3649] <= 1'h0;
      write_enable_data_log_force[3650] <= 1'h0;
      write_enable_data_log_force[3651] <= 1'h0;
      write_enable_data_log_force[3652] <= 1'h0;
      write_enable_data_log_force[3653] <= 1'h0;
      write_enable_data_log_force[3654] <= 1'h0;
      write_enable_data_log_force[3655] <= 1'h0;
      write_enable_data_log_force[3656] <= 1'h0;
      write_enable_data_log_force[3657] <= 1'h0;
      write_enable_data_log_force[3658] <= 1'h0;
      write_enable_data_log_force[3659] <= 1'h0;
      write_enable_data_log_force[3660] <= 1'h0;
      write_enable_data_log_force[3661] <= 1'h0;
      write_enable_data_log_force[3662] <= 1'h0;
      write_enable_data_log_force[3663] <= 1'h0;
      write_enable_data_log_force[3664] <= 1'h0;
      write_enable_data_log_force[3665] <= 1'h0;
      write_enable_data_log_force[3666] <= 1'h0;
      write_enable_data_log_force[3667] <= 1'h0;
      write_enable_data_log_force[3668] <= 1'h0;
      write_enable_data_log_force[3669] <= 1'h0;
      write_enable_data_log_force[3670] <= 1'h0;
      write_enable_data_log_force[3671] <= 1'h0;
      write_enable_data_log_force[3672] <= 1'h0;
      write_enable_data_log_force[3673] <= 1'h0;
      write_enable_data_log_force[3674] <= 1'h0;
      write_enable_data_log_force[3675] <= 1'h0;
      write_enable_data_log_force[3676] <= 1'h0;
      write_enable_data_log_force[3677] <= 1'h0;
      write_enable_data_log_force[3678] <= 1'h0;
      write_enable_data_log_force[3679] <= 1'h0;
      write_enable_data_log_force[3680] <= 1'h0;
      write_enable_data_log_force[3681] <= 1'h0;
      write_enable_data_log_force[3682] <= 1'h0;
      write_enable_data_log_force[3683] <= 1'h0;
      write_enable_data_log_force[3684] <= 1'h0;
      write_enable_data_log_force[3685] <= 1'h0;
      write_enable_data_log_force[3686] <= 1'h0;
      write_enable_data_log_force[3687] <= 1'h0;
      write_enable_data_log_force[3688] <= 1'h0;
      write_enable_data_log_force[3689] <= 1'h0;
      write_enable_data_log_force[3690] <= 1'h0;
      write_enable_data_log_force[3691] <= 1'h0;
      write_enable_data_log_force[3692] <= 1'h0;
      write_enable_data_log_force[3693] <= 1'h0;
      write_enable_data_log_force[3694] <= 1'h0;
      write_enable_data_log_force[3695] <= 1'h0;
      write_enable_data_log_force[3696] <= 1'h0;
      write_enable_data_log_force[3697] <= 1'h0;
      write_enable_data_log_force[3698] <= 1'h0;
      write_enable_data_log_force[3699] <= 1'h0;
      write_enable_data_log_force[3700] <= 1'h0;
      write_enable_data_log_force[3701] <= 1'h0;
      write_enable_data_log_force[3702] <= 1'h0;
      write_enable_data_log_force[3703] <= 1'h0;
      write_enable_data_log_force[3704] <= 1'h0;
      write_enable_data_log_force[3705] <= 1'h0;
      write_enable_data_log_force[3706] <= 1'h0;
      write_enable_data_log_force[3707] <= 1'h0;
      write_enable_data_log_force[3708] <= 1'h0;
      write_enable_data_log_force[3709] <= 1'h0;
      write_enable_data_log_force[3710] <= 1'h0;
      write_enable_data_log_force[3711] <= 1'h0;
      write_enable_data_log_force[3712] <= 1'h0;
      write_enable_data_log_force[3713] <= 1'h0;
      write_enable_data_log_force[3714] <= 1'h0;
      write_enable_data_log_force[3715] <= 1'h0;
      write_enable_data_log_force[3716] <= 1'h0;
      write_enable_data_log_force[3717] <= 1'h0;
      write_enable_data_log_force[3718] <= 1'h0;
      write_enable_data_log_force[3719] <= 1'h0;
      write_enable_data_log_force[3720] <= 1'h0;
      write_enable_data_log_force[3721] <= 1'h0;
      write_enable_data_log_force[3722] <= 1'h0;
      write_enable_data_log_force[3723] <= 1'h0;
      write_enable_data_log_force[3724] <= 1'h0;
      write_enable_data_log_force[3725] <= 1'h0;
      write_enable_data_log_force[3726] <= 1'h0;
      write_enable_data_log_force[3727] <= 1'h0;
      write_enable_data_log_force[3728] <= 1'h0;
      write_enable_data_log_force[3729] <= 1'h0;
      write_enable_data_log_force[3730] <= 1'h0;
      write_enable_data_log_force[3731] <= 1'h0;
      write_enable_data_log_force[3732] <= 1'h0;
      write_enable_data_log_force[3733] <= 1'h0;
      write_enable_data_log_force[3734] <= 1'h0;
      write_enable_data_log_force[3735] <= 1'h0;
      write_enable_data_log_force[3736] <= 1'h0;
      write_enable_data_log_force[3737] <= 1'h0;
      write_enable_data_log_force[3738] <= 1'h0;
      write_enable_data_log_force[3739] <= 1'h0;
      write_enable_data_log_force[3740] <= 1'h0;
      write_enable_data_log_force[3741] <= 1'h0;
      write_enable_data_log_force[3742] <= 1'h0;
      write_enable_data_log_force[3743] <= 1'h0;
      write_enable_data_log_force[3744] <= 1'h0;
      write_enable_data_log_force[3745] <= 1'h0;
      write_enable_data_log_force[3746] <= 1'h0;
      write_enable_data_log_force[3747] <= 1'h0;
      write_enable_data_log_force[3748] <= 1'h0;
      write_enable_data_log_force[3749] <= 1'h0;
      write_enable_data_log_force[3750] <= 1'h0;
      write_enable_data_log_force[3751] <= 1'h0;
      write_enable_data_log_force[3752] <= 1'h0;
      write_enable_data_log_force[3753] <= 1'h0;
      write_enable_data_log_force[3754] <= 1'h0;
      write_enable_data_log_force[3755] <= 1'h0;
      write_enable_data_log_force[3756] <= 1'h0;
      write_enable_data_log_force[3757] <= 1'h0;
      write_enable_data_log_force[3758] <= 1'h0;
      write_enable_data_log_force[3759] <= 1'h0;
      write_enable_data_log_force[3760] <= 1'h0;
      write_enable_data_log_force[3761] <= 1'h0;
      write_enable_data_log_force[3762] <= 1'h0;
      write_enable_data_log_force[3763] <= 1'h0;
      write_enable_data_log_force[3764] <= 1'h0;
      write_enable_data_log_force[3765] <= 1'h0;
      write_enable_data_log_force[3766] <= 1'h0;
      write_enable_data_log_force[3767] <= 1'h0;
      write_enable_data_log_force[3768] <= 1'h0;
      write_enable_data_log_force[3769] <= 1'h0;
      write_enable_data_log_force[3770] <= 1'h0;
      write_enable_data_log_force[3771] <= 1'h0;
      write_enable_data_log_force[3772] <= 1'h0;
      write_enable_data_log_force[3773] <= 1'h0;
      write_enable_data_log_force[3774] <= 1'h0;
      write_enable_data_log_force[3775] <= 1'h0;
      write_enable_data_log_force[3776] <= 1'h0;
      write_enable_data_log_force[3777] <= 1'h0;
      write_enable_data_log_force[3778] <= 1'h0;
      write_enable_data_log_force[3779] <= 1'h0;
      write_enable_data_log_force[3780] <= 1'h0;
      write_enable_data_log_force[3781] <= 1'h0;
      write_enable_data_log_force[3782] <= 1'h0;
      write_enable_data_log_force[3783] <= 1'h0;
      write_enable_data_log_force[3784] <= 1'h0;
      write_enable_data_log_force[3785] <= 1'h0;
      write_enable_data_log_force[3786] <= 1'h0;
      write_enable_data_log_force[3787] <= 1'h0;
      write_enable_data_log_force[3788] <= 1'h0;
      write_enable_data_log_force[3789] <= 1'h0;
      write_enable_data_log_force[3790] <= 1'h0;
      write_enable_data_log_force[3791] <= 1'h0;
      write_enable_data_log_force[3792] <= 1'h0;
      write_enable_data_log_force[3793] <= 1'h0;
      write_enable_data_log_force[3794] <= 1'h0;
      write_enable_data_log_force[3795] <= 1'h0;
      write_enable_data_log_force[3796] <= 1'h0;
      write_enable_data_log_force[3797] <= 1'h0;
      write_enable_data_log_force[3798] <= 1'h0;
      write_enable_data_log_force[3799] <= 1'h0;
      write_enable_data_log_force[3800] <= 1'h0;
      write_enable_data_log_force[3801] <= 1'h0;
      write_enable_data_log_force[3802] <= 1'h0;
      write_enable_data_log_force[3803] <= 1'h0;
      write_enable_data_log_force[3804] <= 1'h0;
      write_enable_data_log_force[3805] <= 1'h0;
      write_enable_data_log_force[3806] <= 1'h0;
      write_enable_data_log_force[3807] <= 1'h0;
      write_enable_data_log_force[3808] <= 1'h0;
      write_enable_data_log_force[3809] <= 1'h0;
      write_enable_data_log_force[3810] <= 1'h0;
      write_enable_data_log_force[3811] <= 1'h0;
      write_enable_data_log_force[3812] <= 1'h0;
      write_enable_data_log_force[3813] <= 1'h0;
      write_enable_data_log_force[3814] <= 1'h0;
      write_enable_data_log_force[3815] <= 1'h0;
      write_enable_data_log_force[3816] <= 1'h0;
      write_enable_data_log_force[3817] <= 1'h0;
      write_enable_data_log_force[3818] <= 1'h0;
      write_enable_data_log_force[3819] <= 1'h0;
      write_enable_data_log_force[3820] <= 1'h0;
      write_enable_data_log_force[3821] <= 1'h0;
      write_enable_data_log_force[3822] <= 1'h0;
      write_enable_data_log_force[3823] <= 1'h0;
      write_enable_data_log_force[3824] <= 1'h0;
      write_enable_data_log_force[3825] <= 1'h0;
      write_enable_data_log_force[3826] <= 1'h0;
      write_enable_data_log_force[3827] <= 1'h0;
      write_enable_data_log_force[3828] <= 1'h0;
      write_enable_data_log_force[3829] <= 1'h0;
      write_enable_data_log_force[3830] <= 1'h0;
      write_enable_data_log_force[3831] <= 1'h0;
      write_enable_data_log_force[3832] <= 1'h0;
      write_enable_data_log_force[3833] <= 1'h0;
      write_enable_data_log_force[3834] <= 1'h0;
      write_enable_data_log_force[3835] <= 1'h0;
      write_enable_data_log_force[3836] <= 1'h0;
      write_enable_data_log_force[3837] <= 1'h0;
      write_enable_data_log_force[3838] <= 1'h0;
      write_enable_data_log_force[3839] <= 1'h0;
      write_enable_data_log_force[3840] <= 1'h0;
      write_enable_data_log_force[3841] <= 1'h0;
      write_enable_data_log_force[3842] <= 1'h0;
      write_enable_data_log_force[3843] <= 1'h0;
      write_enable_data_log_force[3844] <= 1'h0;
      write_enable_data_log_force[3845] <= 1'h0;
      write_enable_data_log_force[3846] <= 1'h0;
      write_enable_data_log_force[3847] <= 1'h0;
      write_enable_data_log_force[3848] <= 1'h0;
      write_enable_data_log_force[3849] <= 1'h0;
      write_enable_data_log_force[3850] <= 1'h0;
      write_enable_data_log_force[3851] <= 1'h0;
      write_enable_data_log_force[3852] <= 1'h0;
      write_enable_data_log_force[3853] <= 1'h0;
      write_enable_data_log_force[3854] <= 1'h0;
      write_enable_data_log_force[3855] <= 1'h0;
      write_enable_data_log_force[3856] <= 1'h0;
      write_enable_data_log_force[3857] <= 1'h0;
      write_enable_data_log_force[3858] <= 1'h0;
      write_enable_data_log_force[3859] <= 1'h0;
      write_enable_data_log_force[3860] <= 1'h0;
      write_enable_data_log_force[3861] <= 1'h0;
      write_enable_data_log_force[3862] <= 1'h0;
      write_enable_data_log_force[3863] <= 1'h0;
      write_enable_data_log_force[3864] <= 1'h0;
      write_enable_data_log_force[3865] <= 1'h0;
      write_enable_data_log_force[3866] <= 1'h0;
      write_enable_data_log_force[3867] <= 1'h0;
      write_enable_data_log_force[3868] <= 1'h0;
      write_enable_data_log_force[3869] <= 1'h0;
      write_enable_data_log_force[3870] <= 1'h0;
      write_enable_data_log_force[3871] <= 1'h0;
      write_enable_data_log_force[3872] <= 1'h0;
      write_enable_data_log_force[3873] <= 1'h0;
      write_enable_data_log_force[3874] <= 1'h0;
      write_enable_data_log_force[3875] <= 1'h0;
      write_enable_data_log_force[3876] <= 1'h0;
      write_enable_data_log_force[3877] <= 1'h0;
      write_enable_data_log_force[3878] <= 1'h0;
      write_enable_data_log_force[3879] <= 1'h0;
      write_enable_data_log_force[3880] <= 1'h0;
      write_enable_data_log_force[3881] <= 1'h0;
      write_enable_data_log_force[3882] <= 1'h0;
      write_enable_data_log_force[3883] <= 1'h0;
      write_enable_data_log_force[3884] <= 1'h0;
      write_enable_data_log_force[3885] <= 1'h0;
      write_enable_data_log_force[3886] <= 1'h0;
      write_enable_data_log_force[3887] <= 1'h0;
      write_enable_data_log_force[3888] <= 1'h0;
      write_enable_data_log_force[3889] <= 1'h0;
      write_enable_data_log_force[3890] <= 1'h0;
      write_enable_data_log_force[3891] <= 1'h0;
      write_enable_data_log_force[3892] <= 1'h0;
      write_enable_data_log_force[3893] <= 1'h0;
      write_enable_data_log_force[3894] <= 1'h0;
      write_enable_data_log_force[3895] <= 1'h0;
      write_enable_data_log_force[3896] <= 1'h0;
      write_enable_data_log_force[3897] <= 1'h0;
      write_enable_data_log_force[3898] <= 1'h0;
      write_enable_data_log_force[3899] <= 1'h0;
      write_enable_data_log_force[3900] <= 1'h0;
      write_enable_data_log_force[3901] <= 1'h0;
      write_enable_data_log_force[3902] <= 1'h0;
      write_enable_data_log_force[3903] <= 1'h0;
      write_enable_data_log_force[3904] <= 1'h0;
      write_enable_data_log_force[3905] <= 1'h0;
      write_enable_data_log_force[3906] <= 1'h0;
      write_enable_data_log_force[3907] <= 1'h0;
      write_enable_data_log_force[3908] <= 1'h0;
      write_enable_data_log_force[3909] <= 1'h0;
      write_enable_data_log_force[3910] <= 1'h0;
      write_enable_data_log_force[3911] <= 1'h0;
      write_enable_data_log_force[3912] <= 1'h0;
      write_enable_data_log_force[3913] <= 1'h0;
      write_enable_data_log_force[3914] <= 1'h0;
      write_enable_data_log_force[3915] <= 1'h0;
      write_enable_data_log_force[3916] <= 1'h0;
      write_enable_data_log_force[3917] <= 1'h0;
      write_enable_data_log_force[3918] <= 1'h0;
      write_enable_data_log_force[3919] <= 1'h0;
      write_enable_data_log_force[3920] <= 1'h0;
      write_enable_data_log_force[3921] <= 1'h0;
      write_enable_data_log_force[3922] <= 1'h0;
      write_enable_data_log_force[3923] <= 1'h0;
      write_enable_data_log_force[3924] <= 1'h0;
      write_enable_data_log_force[3925] <= 1'h0;
      write_enable_data_log_force[3926] <= 1'h0;
      write_enable_data_log_force[3927] <= 1'h0;
      write_enable_data_log_force[3928] <= 1'h0;
      write_enable_data_log_force[3929] <= 1'h0;
      write_enable_data_log_force[3930] <= 1'h0;
      write_enable_data_log_force[3931] <= 1'h0;
      write_enable_data_log_force[3932] <= 1'h0;
      write_enable_data_log_force[3933] <= 1'h0;
      write_enable_data_log_force[3934] <= 1'h0;
      write_enable_data_log_force[3935] <= 1'h0;
      write_enable_data_log_force[3936] <= 1'h0;
      write_enable_data_log_force[3937] <= 1'h0;
      write_enable_data_log_force[3938] <= 1'h0;
      write_enable_data_log_force[3939] <= 1'h0;
      write_enable_data_log_force[3940] <= 1'h0;
      write_enable_data_log_force[3941] <= 1'h0;
      write_enable_data_log_force[3942] <= 1'h0;
      write_enable_data_log_force[3943] <= 1'h0;
      write_enable_data_log_force[3944] <= 1'h0;
      write_enable_data_log_force[3945] <= 1'h0;
      write_enable_data_log_force[3946] <= 1'h0;
      write_enable_data_log_force[3947] <= 1'h0;
      write_enable_data_log_force[3948] <= 1'h0;
      write_enable_data_log_force[3949] <= 1'h0;
      write_enable_data_log_force[3950] <= 1'h0;
      write_enable_data_log_force[3951] <= 1'h0;
      write_enable_data_log_force[3952] <= 1'h0;
      write_enable_data_log_force[3953] <= 1'h0;
      write_enable_data_log_force[3954] <= 1'h0;
      write_enable_data_log_force[3955] <= 1'h0;
      write_enable_data_log_force[3956] <= 1'h0;
      write_enable_data_log_force[3957] <= 1'h0;
      write_enable_data_log_force[3958] <= 1'h0;
      write_enable_data_log_force[3959] <= 1'h0;
      write_enable_data_log_force[3960] <= 1'h0;
      write_enable_data_log_force[3961] <= 1'h0;
      write_enable_data_log_force[3962] <= 1'h0;
      write_enable_data_log_force[3963] <= 1'h0;
      write_enable_data_log_force[3964] <= 1'h0;
      write_enable_data_log_force[3965] <= 1'h0;
      write_enable_data_log_force[3966] <= 1'h0;
      write_enable_data_log_force[3967] <= 1'h0;
      write_enable_data_log_force[3968] <= 1'h0;
      write_enable_data_log_force[3969] <= 1'h0;
      write_enable_data_log_force[3970] <= 1'h0;
      write_enable_data_log_force[3971] <= 1'h0;
      write_enable_data_log_force[3972] <= 1'h0;
      write_enable_data_log_force[3973] <= 1'h0;
      write_enable_data_log_force[3974] <= 1'h0;
      write_enable_data_log_force[3975] <= 1'h0;
      write_enable_data_log_force[3976] <= 1'h0;
      write_enable_data_log_force[3977] <= 1'h0;
      write_enable_data_log_force[3978] <= 1'h0;
      write_enable_data_log_force[3979] <= 1'h0;
      write_enable_data_log_force[3980] <= 1'h0;
      write_enable_data_log_force[3981] <= 1'h0;
      write_enable_data_log_force[3982] <= 1'h0;
      write_enable_data_log_force[3983] <= 1'h0;
      write_enable_data_log_force[3984] <= 1'h0;
      write_enable_data_log_force[3985] <= 1'h0;
      write_enable_data_log_force[3986] <= 1'h0;
      write_enable_data_log_force[3987] <= 1'h0;
      write_enable_data_log_force[3988] <= 1'h0;
      write_enable_data_log_force[3989] <= 1'h0;
      write_enable_data_log_force[3990] <= 1'h0;
      write_enable_data_log_force[3991] <= 1'h0;
      write_enable_data_log_force[3992] <= 1'h0;
      write_enable_data_log_force[3993] <= 1'h0;
      write_enable_data_log_force[3994] <= 1'h0;
      write_enable_data_log_force[3995] <= 1'h0;
      write_enable_data_log_force[3996] <= 1'h0;
      write_enable_data_log_force[3997] <= 1'h0;
      write_enable_data_log_force[3998] <= 1'h0;
      write_enable_data_log_force[3999] <= 1'h0;
      write_enable_data_log_force[4000] <= 1'h0;
      write_enable_data_log_force[4001] <= 1'h0;
      write_enable_data_log_force[4002] <= 1'h0;
      write_enable_data_log_force[4003] <= 1'h0;
      write_enable_data_log_force[4004] <= 1'h0;
      write_enable_data_log_force[4005] <= 1'h0;
      write_enable_data_log_force[4006] <= 1'h0;
      write_enable_data_log_force[4007] <= 1'h0;
      write_enable_data_log_force[4008] <= 1'h0;
      write_enable_data_log_force[4009] <= 1'h0;
      write_enable_data_log_force[4010] <= 1'h0;
      write_enable_data_log_force[4011] <= 1'h0;
      write_enable_data_log_force[4012] <= 1'h0;
      write_enable_data_log_force[4013] <= 1'h0;
      write_enable_data_log_force[4014] <= 1'h0;
      write_enable_data_log_force[4015] <= 1'h0;
      write_enable_data_log_force[4016] <= 1'h0;
      write_enable_data_log_force[4017] <= 1'h0;
      write_enable_data_log_force[4018] <= 1'h0;
      write_enable_data_log_force[4019] <= 1'h0;
      write_enable_data_log_force[4020] <= 1'h0;
      write_enable_data_log_force[4021] <= 1'h0;
      write_enable_data_log_force[4022] <= 1'h0;
      write_enable_data_log_force[4023] <= 1'h0;
      write_enable_data_log_force[4024] <= 1'h0;
      write_enable_data_log_force[4025] <= 1'h0;
      write_enable_data_log_force[4026] <= 1'h0;
      write_enable_data_log_force[4027] <= 1'h0;
      write_enable_data_log_force[4028] <= 1'h0;
      write_enable_data_log_force[4029] <= 1'h0;
      write_enable_data_log_force[4030] <= 1'h0;
      write_enable_data_log_force[4031] <= 1'h0;
      write_enable_data_log_force[4032] <= 1'h0;
      write_enable_data_log_force[4033] <= 1'h0;
      write_enable_data_log_force[4034] <= 1'h0;
      write_enable_data_log_force[4035] <= 1'h0;
      write_enable_data_log_force[4036] <= 1'h0;
      write_enable_data_log_force[4037] <= 1'h0;
      write_enable_data_log_force[4038] <= 1'h0;
      write_enable_data_log_force[4039] <= 1'h0;
      write_enable_data_log_force[4040] <= 1'h0;
      write_enable_data_log_force[4041] <= 1'h0;
      write_enable_data_log_force[4042] <= 1'h0;
      write_enable_data_log_force[4043] <= 1'h0;
      write_enable_data_log_force[4044] <= 1'h0;
      write_enable_data_log_force[4045] <= 1'h0;
      write_enable_data_log_force[4046] <= 1'h0;
      write_enable_data_log_force[4047] <= 1'h0;
      write_enable_data_log_force[4048] <= 1'h0;
      write_enable_data_log_force[4049] <= 1'h0;
      write_enable_data_log_force[4050] <= 1'h0;
      write_enable_data_log_force[4051] <= 1'h0;
      write_enable_data_log_force[4052] <= 1'h0;
      write_enable_data_log_force[4053] <= 1'h0;
      write_enable_data_log_force[4054] <= 1'h0;
      write_enable_data_log_force[4055] <= 1'h0;
      write_enable_data_log_force[4056] <= 1'h0;
      write_enable_data_log_force[4057] <= 1'h0;
      write_enable_data_log_force[4058] <= 1'h0;
      write_enable_data_log_force[4059] <= 1'h0;
      write_enable_data_log_force[4060] <= 1'h0;
      write_enable_data_log_force[4061] <= 1'h0;
      write_enable_data_log_force[4062] <= 1'h0;
      write_enable_data_log_force[4063] <= 1'h0;
      write_enable_data_log_force[4064] <= 1'h0;
      write_enable_data_log_force[4065] <= 1'h0;
      write_enable_data_log_force[4066] <= 1'h0;
      write_enable_data_log_force[4067] <= 1'h0;
      write_enable_data_log_force[4068] <= 1'h0;
      write_enable_data_log_force[4069] <= 1'h0;
      write_enable_data_log_force[4070] <= 1'h0;
      write_enable_data_log_force[4071] <= 1'h0;
      write_enable_data_log_force[4072] <= 1'h0;
      write_enable_data_log_force[4073] <= 1'h0;
      write_enable_data_log_force[4074] <= 1'h0;
      write_enable_data_log_force[4075] <= 1'h0;
      write_enable_data_log_force[4076] <= 1'h0;
      write_enable_data_log_force[4077] <= 1'h0;
      write_enable_data_log_force[4078] <= 1'h0;
      write_enable_data_log_force[4079] <= 1'h0;
      write_enable_data_log_force[4080] <= 1'h0;
      write_enable_data_log_force[4081] <= 1'h0;
      write_enable_data_log_force[4082] <= 1'h0;
      write_enable_data_log_force[4083] <= 1'h0;
      write_enable_data_log_force[4084] <= 1'h0;
      write_enable_data_log_force[4085] <= 1'h0;
      write_enable_data_log_force[4086] <= 1'h0;
      write_enable_data_log_force[4087] <= 1'h0;
      write_enable_data_log_force[4088] <= 1'h0;
      write_enable_data_log_force[4089] <= 1'h0;
      write_enable_data_log_force[4090] <= 1'h0;
      write_enable_data_log_force[4091] <= 1'h0;
      write_enable_data_log_force[4092] <= 1'h0;
      write_enable_data_log_force[4093] <= 1'h0;
      write_enable_data_log_force[4094] <= 1'h0;
      write_enable_data_log_force[4095] <= 1'h0;
      write_enable_data_log_force[4096] <= 1'h0;
      write_enable_data_log_force[4097] <= 1'h0;
      write_enable_data_log_force[4098] <= 1'h0;
      write_enable_data_log_force[4099] <= 1'h0;
      write_enable_data_log_force[4100] <= 1'h0;
      write_enable_data_log_force[4101] <= 1'h0;
      write_enable_data_log_force[4102] <= 1'h0;
      write_enable_data_log_force[4103] <= 1'h0;
      write_enable_data_log_force[4104] <= 1'h0;
      write_enable_data_log_force[4105] <= 1'h0;
      write_enable_data_log_force[4106] <= 1'h0;
      write_enable_data_log_force[4107] <= 1'h0;
      write_enable_data_log_force[4108] <= 1'h0;
      write_enable_data_log_force[4109] <= 1'h0;
      write_enable_data_log_force[4110] <= 1'h0;
      write_enable_data_log_force[4111] <= 1'h0;
      write_enable_data_log_force[4112] <= 1'h0;
      write_enable_data_log_force[4113] <= 1'h0;
      write_enable_data_log_force[4114] <= 1'h0;
      write_enable_data_log_force[4115] <= 1'h0;
      write_enable_data_log_force[4116] <= 1'h0;
      write_enable_data_log_force[4117] <= 1'h0;
      write_enable_data_log_force[4118] <= 1'h0;
      write_enable_data_log_force[4119] <= 1'h0;
      write_enable_data_log_force[4120] <= 1'h0;
      write_enable_data_log_force[4121] <= 1'h0;
      write_enable_data_log_force[4122] <= 1'h0;
      write_enable_data_log_force[4123] <= 1'h0;
      write_enable_data_log_force[4124] <= 1'h0;
      write_enable_data_log_force[4125] <= 1'h0;
      write_enable_data_log_force[4126] <= 1'h0;
      write_enable_data_log_force[4127] <= 1'h0;
      write_enable_data_log_force[4128] <= 1'h0;
      write_enable_data_log_force[4129] <= 1'h0;
      write_enable_data_log_force[4130] <= 1'h0;
      write_enable_data_log_force[4131] <= 1'h0;
      write_enable_data_log_force[4132] <= 1'h0;
      write_enable_data_log_force[4133] <= 1'h0;
      write_enable_data_log_force[4134] <= 1'h0;
      write_enable_data_log_force[4135] <= 1'h0;
      write_enable_data_log_force[4136] <= 1'h0;
      write_enable_data_log_force[4137] <= 1'h0;
      write_enable_data_log_force[4138] <= 1'h0;
      write_enable_data_log_force[4139] <= 1'h0;
      write_enable_data_log_force[4140] <= 1'h0;
      write_enable_data_log_force[4141] <= 1'h0;
      write_enable_data_log_force[4142] <= 1'h0;
      write_enable_data_log_force[4143] <= 1'h0;
      write_enable_data_log_force[4144] <= 1'h0;
      write_enable_data_log_force[4145] <= 1'h0;
      write_enable_data_log_force[4146] <= 1'h0;
      write_enable_data_log_force[4147] <= 1'h0;
      write_enable_data_log_force[4148] <= 1'h0;
      write_enable_data_log_force[4149] <= 1'h0;
      write_enable_data_log_force[4150] <= 1'h0;
      write_enable_data_log_force[4151] <= 1'h0;
      write_enable_data_log_force[4152] <= 1'h0;
      write_enable_data_log_force[4153] <= 1'h0;
      write_enable_data_log_force[4154] <= 1'h0;
      write_enable_data_log_force[4155] <= 1'h0;
      write_enable_data_log_force[4156] <= 1'h0;
      write_enable_data_log_force[4157] <= 1'h0;
      write_enable_data_log_force[4158] <= 1'h0;
      write_enable_data_log_force[4159] <= 1'h0;
      write_enable_data_log_force[4160] <= 1'h0;
      write_enable_data_log_force[4161] <= 1'h0;
      write_enable_data_log_force[4162] <= 1'h0;
      write_enable_data_log_force[4163] <= 1'h0;
      write_enable_data_log_force[4164] <= 1'h0;
      write_enable_data_log_force[4165] <= 1'h0;
      write_enable_data_log_force[4166] <= 1'h0;
      write_enable_data_log_force[4167] <= 1'h0;
      write_enable_data_log_force[4168] <= 1'h0;
      write_enable_data_log_force[4169] <= 1'h0;
      write_enable_data_log_force[4170] <= 1'h0;
      write_enable_data_log_force[4171] <= 1'h0;
      write_enable_data_log_force[4172] <= 1'h0;
      write_enable_data_log_force[4173] <= 1'h0;
      write_enable_data_log_force[4174] <= 1'h0;
      write_enable_data_log_force[4175] <= 1'h0;
      write_enable_data_log_force[4176] <= 1'h0;
      write_enable_data_log_force[4177] <= 1'h0;
      write_enable_data_log_force[4178] <= 1'h0;
      write_enable_data_log_force[4179] <= 1'h0;
      write_enable_data_log_force[4180] <= 1'h0;
      write_enable_data_log_force[4181] <= 1'h0;
      write_enable_data_log_force[4182] <= 1'h0;
      write_enable_data_log_force[4183] <= 1'h0;
      write_enable_data_log_force[4184] <= 1'h0;
      write_enable_data_log_force[4185] <= 1'h0;
      write_enable_data_log_force[4186] <= 1'h0;
      write_enable_data_log_force[4187] <= 1'h0;
      write_enable_data_log_force[4188] <= 1'h0;
      write_enable_data_log_force[4189] <= 1'h0;
      write_enable_data_log_force[4190] <= 1'h0;
      write_enable_data_log_force[4191] <= 1'h0;
      write_enable_data_log_force[4192] <= 1'h0;
      write_enable_data_log_force[4193] <= 1'h0;
      write_enable_data_log_force[4194] <= 1'h0;
      write_enable_data_log_force[4195] <= 1'h0;
      write_enable_data_log_force[4196] <= 1'h0;
      write_enable_data_log_force[4197] <= 1'h0;
      write_enable_data_log_force[4198] <= 1'h0;
      write_enable_data_log_force[4199] <= 1'h0;
      write_enable_data_log_force[4200] <= 1'h0;
      write_enable_data_log_force[4201] <= 1'h0;
      write_enable_data_log_force[4202] <= 1'h0;
      write_enable_data_log_force[4203] <= 1'h0;
      write_enable_data_log_force[4204] <= 1'h0;
      write_enable_data_log_force[4205] <= 1'h0;
      write_enable_data_log_force[4206] <= 1'h0;
      write_enable_data_log_force[4207] <= 1'h0;
      write_enable_data_log_force[4208] <= 1'h0;
      write_enable_data_log_force[4209] <= 1'h0;
      write_enable_data_log_force[4210] <= 1'h0;
      write_enable_data_log_force[4211] <= 1'h0;
      write_enable_data_log_force[4212] <= 1'h0;
      write_enable_data_log_force[4213] <= 1'h0;
      write_enable_data_log_force[4214] <= 1'h0;
      write_enable_data_log_force[4215] <= 1'h0;
      write_enable_data_log_force[4216] <= 1'h0;
      write_enable_data_log_force[4217] <= 1'h0;
      write_enable_data_log_force[4218] <= 1'h0;
      write_enable_data_log_force[4219] <= 1'h0;
      write_enable_data_log_force[4220] <= 1'h0;
      write_enable_data_log_force[4221] <= 1'h0;
      write_enable_data_log_force[4222] <= 1'h0;
      write_enable_data_log_force[4223] <= 1'h0;
      write_enable_data_log_force[4224] <= 1'h0;
      write_enable_data_log_force[4225] <= 1'h0;
      write_enable_data_log_force[4226] <= 1'h0;
      write_enable_data_log_force[4227] <= 1'h0;
      write_enable_data_log_force[4228] <= 1'h0;
      write_enable_data_log_force[4229] <= 1'h0;
      write_enable_data_log_force[4230] <= 1'h0;
      write_enable_data_log_force[4231] <= 1'h0;
      write_enable_data_log_force[4232] <= 1'h0;
      write_enable_data_log_force[4233] <= 1'h0;
      write_enable_data_log_force[4234] <= 1'h0;
      write_enable_data_log_force[4235] <= 1'h0;
      write_enable_data_log_force[4236] <= 1'h0;
      write_enable_data_log_force[4237] <= 1'h0;
      write_enable_data_log_force[4238] <= 1'h0;
      write_enable_data_log_force[4239] <= 1'h0;
      write_enable_data_log_force[4240] <= 1'h0;
      write_enable_data_log_force[4241] <= 1'h0;
      write_enable_data_log_force[4242] <= 1'h0;
      write_enable_data_log_force[4243] <= 1'h0;
      write_enable_data_log_force[4244] <= 1'h0;
      write_enable_data_log_force[4245] <= 1'h0;
      write_enable_data_log_force[4246] <= 1'h0;
      write_enable_data_log_force[4247] <= 1'h0;
      write_enable_data_log_force[4248] <= 1'h0;
      write_enable_data_log_force[4249] <= 1'h0;
      write_enable_data_log_force[4250] <= 1'h0;
      write_enable_data_log_force[4251] <= 1'h0;
      write_enable_data_log_force[4252] <= 1'h0;
      write_enable_data_log_force[4253] <= 1'h0;
      write_enable_data_log_force[4254] <= 1'h0;
      write_enable_data_log_force[4255] <= 1'h0;
      write_enable_data_log_force[4256] <= 1'h0;
      write_enable_data_log_force[4257] <= 1'h0;
      write_enable_data_log_force[4258] <= 1'h0;
      write_enable_data_log_force[4259] <= 1'h0;
      write_enable_data_log_force[4260] <= 1'h0;
      write_enable_data_log_force[4261] <= 1'h0;
      write_enable_data_log_force[4262] <= 1'h0;
      write_enable_data_log_force[4263] <= 1'h0;
      write_enable_data_log_force[4264] <= 1'h0;
      write_enable_data_log_force[4265] <= 1'h0;
      write_enable_data_log_force[4266] <= 1'h0;
      write_enable_data_log_force[4267] <= 1'h0;
      write_enable_data_log_force[4268] <= 1'h0;
      write_enable_data_log_force[4269] <= 1'h0;
      write_enable_data_log_force[4270] <= 1'h0;
      write_enable_data_log_force[4271] <= 1'h0;
      write_enable_data_log_force[4272] <= 1'h0;
      write_enable_data_log_force[4273] <= 1'h0;
      write_enable_data_log_force[4274] <= 1'h0;
      write_enable_data_log_force[4275] <= 1'h0;
      write_enable_data_log_force[4276] <= 1'h0;
      write_enable_data_log_force[4277] <= 1'h0;
      write_enable_data_log_force[4278] <= 1'h0;
      write_enable_data_log_force[4279] <= 1'h0;
      write_enable_data_log_force[4280] <= 1'h0;
      write_enable_data_log_force[4281] <= 1'h0;
      write_enable_data_log_force[4282] <= 1'h0;
      write_enable_data_log_force[4283] <= 1'h0;
      write_enable_data_log_force[4284] <= 1'h0;
      write_enable_data_log_force[4285] <= 1'h0;
      write_enable_data_log_force[4286] <= 1'h0;
      write_enable_data_log_force[4287] <= 1'h0;
      write_enable_data_log_force[4288] <= 1'h0;
      write_enable_data_log_force[4289] <= 1'h0;
      write_enable_data_log_force[4290] <= 1'h0;
      write_enable_data_log_force[4291] <= 1'h0;
      write_enable_data_log_force[4292] <= 1'h0;
      write_enable_data_log_force[4293] <= 1'h0;
      write_enable_data_log_force[4294] <= 1'h0;
      write_enable_data_log_force[4295] <= 1'h0;
      write_enable_data_log_force[4296] <= 1'h0;
      write_enable_data_log_force[4297] <= 1'h0;
      write_enable_data_log_force[4298] <= 1'h0;
      write_enable_data_log_force[4299] <= 1'h0;
      write_enable_data_log_force[4300] <= 1'h0;
      write_enable_data_log_force[4301] <= 1'h0;
      write_enable_data_log_force[4302] <= 1'h0;
      write_enable_data_log_force[4303] <= 1'h0;
      write_enable_data_log_force[4304] <= 1'h0;
      write_enable_data_log_force[4305] <= 1'h0;
      write_enable_data_log_force[4306] <= 1'h0;
      write_enable_data_log_force[4307] <= 1'h0;
      write_enable_data_log_force[4308] <= 1'h0;
      write_enable_data_log_force[4309] <= 1'h0;
      write_enable_data_log_force[4310] <= 1'h0;
      write_enable_data_log_force[4311] <= 1'h0;
      write_enable_data_log_force[4312] <= 1'h0;
      write_enable_data_log_force[4313] <= 1'h0;
      write_enable_data_log_force[4314] <= 1'h0;
      write_enable_data_log_force[4315] <= 1'h0;
      write_enable_data_log_force[4316] <= 1'h0;
      write_enable_data_log_force[4317] <= 1'h0;
      write_enable_data_log_force[4318] <= 1'h0;
      write_enable_data_log_force[4319] <= 1'h0;
      write_enable_data_log_force[4320] <= 1'h0;
      write_enable_data_log_force[4321] <= 1'h0;
      write_enable_data_log_force[4322] <= 1'h0;
      write_enable_data_log_force[4323] <= 1'h0;
      write_enable_data_log_force[4324] <= 1'h0;
      write_enable_data_log_force[4325] <= 1'h0;
      write_enable_data_log_force[4326] <= 1'h0;
      write_enable_data_log_force[4327] <= 1'h0;
      write_enable_data_log_force[4328] <= 1'h0;
      write_enable_data_log_force[4329] <= 1'h0;
      write_enable_data_log_force[4330] <= 1'h0;
      write_enable_data_log_force[4331] <= 1'h0;
      write_enable_data_log_force[4332] <= 1'h0;
      write_enable_data_log_force[4333] <= 1'h0;
      write_enable_data_log_force[4334] <= 1'h0;
      write_enable_data_log_force[4335] <= 1'h0;
      write_enable_data_log_force[4336] <= 1'h0;
      write_enable_data_log_force[4337] <= 1'h0;
      write_enable_data_log_force[4338] <= 1'h0;
      write_enable_data_log_force[4339] <= 1'h0;
      write_enable_data_log_force[4340] <= 1'h0;
      write_enable_data_log_force[4341] <= 1'h0;
      write_enable_data_log_force[4342] <= 1'h0;
      write_enable_data_log_force[4343] <= 1'h0;
      write_enable_data_log_force[4344] <= 1'h0;
      write_enable_data_log_force[4345] <= 1'h0;
      write_enable_data_log_force[4346] <= 1'h0;
      write_enable_data_log_force[4347] <= 1'h0;
      write_enable_data_log_force[4348] <= 1'h0;
      write_enable_data_log_force[4349] <= 1'h0;
      write_enable_data_log_force[4350] <= 1'h0;
      write_enable_data_log_force[4351] <= 1'h0;
      write_enable_data_log_force[4352] <= 1'h0;
      write_enable_data_log_force[4353] <= 1'h0;
      write_enable_data_log_force[4354] <= 1'h0;
      write_enable_data_log_force[4355] <= 1'h0;
      write_enable_data_log_force[4356] <= 1'h0;
      write_enable_data_log_force[4357] <= 1'h0;
      write_enable_data_log_force[4358] <= 1'h0;
      write_enable_data_log_force[4359] <= 1'h0;
      write_enable_data_log_force[4360] <= 1'h0;
      write_enable_data_log_force[4361] <= 1'h0;
      write_enable_data_log_force[4362] <= 1'h0;
      write_enable_data_log_force[4363] <= 1'h0;
      write_enable_data_log_force[4364] <= 1'h0;
      write_enable_data_log_force[4365] <= 1'h0;
      write_enable_data_log_force[4366] <= 1'h0;
      write_enable_data_log_force[4367] <= 1'h0;
      write_enable_data_log_force[4368] <= 1'h0;
      write_enable_data_log_force[4369] <= 1'h0;
      write_enable_data_log_force[4370] <= 1'h0;
      write_enable_data_log_force[4371] <= 1'h0;
      write_enable_data_log_force[4372] <= 1'h0;
      write_enable_data_log_force[4373] <= 1'h0;
      write_enable_data_log_force[4374] <= 1'h0;
      write_enable_data_log_force[4375] <= 1'h0;
      write_enable_data_log_force[4376] <= 1'h0;
      write_enable_data_log_force[4377] <= 1'h0;
      write_enable_data_log_force[4378] <= 1'h0;
      write_enable_data_log_force[4379] <= 1'h0;
      write_enable_data_log_force[4380] <= 1'h0;
      write_enable_data_log_force[4381] <= 1'h0;
      write_enable_data_log_force[4382] <= 1'h0;
      write_enable_data_log_force[4383] <= 1'h0;
      write_enable_data_log_force[4384] <= 1'h0;
      write_enable_data_log_force[4385] <= 1'h0;
      write_enable_data_log_force[4386] <= 1'h0;
      write_enable_data_log_force[4387] <= 1'h0;
      write_enable_data_log_force[4388] <= 1'h0;
      write_enable_data_log_force[4389] <= 1'h0;
      write_enable_data_log_force[4390] <= 1'h0;
      write_enable_data_log_force[4391] <= 1'h0;
      write_enable_data_log_force[4392] <= 1'h0;
      write_enable_data_log_force[4393] <= 1'h0;
      write_enable_data_log_force[4394] <= 1'h0;
      write_enable_data_log_force[4395] <= 1'h0;
      write_enable_data_log_force[4396] <= 1'h0;
      write_enable_data_log_force[4397] <= 1'h0;
      write_enable_data_log_force[4398] <= 1'h0;
      write_enable_data_log_force[4399] <= 1'h0;
      write_enable_data_log_force[4400] <= 1'h0;
      write_enable_data_log_force[4401] <= 1'h0;
      write_enable_data_log_force[4402] <= 1'h0;
      write_enable_data_log_force[4403] <= 1'h0;
      write_enable_data_log_force[4404] <= 1'h0;
      write_enable_data_log_force[4405] <= 1'h0;
      write_enable_data_log_force[4406] <= 1'h0;
      write_enable_data_log_force[4407] <= 1'h0;
      write_enable_data_log_force[4408] <= 1'h0;
      write_enable_data_log_force[4409] <= 1'h0;
      write_enable_data_log_force[4410] <= 1'h0;
      write_enable_data_log_force[4411] <= 1'h0;
      write_enable_data_log_force[4412] <= 1'h0;
      write_enable_data_log_force[4413] <= 1'h0;
      write_enable_data_log_force[4414] <= 1'h0;
      write_enable_data_log_force[4415] <= 1'h0;
      write_enable_data_log_force[4416] <= 1'h0;
      write_enable_data_log_force[4417] <= 1'h0;
      write_enable_data_log_force[4418] <= 1'h0;
      write_enable_data_log_force[4419] <= 1'h0;
      write_enable_data_log_force[4420] <= 1'h0;
      write_enable_data_log_force[4421] <= 1'h0;
      write_enable_data_log_force[4422] <= 1'h0;
      write_enable_data_log_force[4423] <= 1'h0;
      write_enable_data_log_force[4424] <= 1'h0;
      write_enable_data_log_force[4425] <= 1'h0;
      write_enable_data_log_force[4426] <= 1'h0;
      write_enable_data_log_force[4427] <= 1'h0;
      write_enable_data_log_force[4428] <= 1'h0;
      write_enable_data_log_force[4429] <= 1'h0;
      write_enable_data_log_force[4430] <= 1'h0;
      write_enable_data_log_force[4431] <= 1'h0;
      write_enable_data_log_force[4432] <= 1'h0;
      write_enable_data_log_force[4433] <= 1'h0;
      write_enable_data_log_force[4434] <= 1'h0;
      write_enable_data_log_force[4435] <= 1'h0;
      write_enable_data_log_force[4436] <= 1'h0;
      write_enable_data_log_force[4437] <= 1'h0;
      write_enable_data_log_force[4438] <= 1'h0;
      write_enable_data_log_force[4439] <= 1'h0;
      write_enable_data_log_force[4440] <= 1'h0;
      write_enable_data_log_force[4441] <= 1'h0;
      write_enable_data_log_force[4442] <= 1'h0;
      write_enable_data_log_force[4443] <= 1'h0;
      write_enable_data_log_force[4444] <= 1'h0;
      write_enable_data_log_force[4445] <= 1'h0;
      write_enable_data_log_force[4446] <= 1'h0;
      write_enable_data_log_force[4447] <= 1'h0;
      write_enable_data_log_force[4448] <= 1'h0;
      write_enable_data_log_force[4449] <= 1'h0;
      write_enable_data_log_force[4450] <= 1'h0;
      write_enable_data_log_force[4451] <= 1'h0;
      write_enable_data_log_force[4452] <= 1'h0;
      write_enable_data_log_force[4453] <= 1'h0;
      write_enable_data_log_force[4454] <= 1'h0;
      write_enable_data_log_force[4455] <= 1'h0;
      write_enable_data_log_force[4456] <= 1'h0;
      write_enable_data_log_force[4457] <= 1'h0;
      write_enable_data_log_force[4458] <= 1'h0;
      write_enable_data_log_force[4459] <= 1'h0;
      write_enable_data_log_force[4460] <= 1'h0;
      write_enable_data_log_force[4461] <= 1'h0;
      write_enable_data_log_force[4462] <= 1'h0;
      write_enable_data_log_force[4463] <= 1'h0;
      write_enable_data_log_force[4464] <= 1'h0;
      write_enable_data_log_force[4465] <= 1'h0;
      write_enable_data_log_force[4466] <= 1'h0;
      write_enable_data_log_force[4467] <= 1'h0;
      write_enable_data_log_force[4468] <= 1'h0;
      write_enable_data_log_force[4469] <= 1'h0;
      write_enable_data_log_force[4470] <= 1'h0;
      write_enable_data_log_force[4471] <= 1'h0;
      write_enable_data_log_force[4472] <= 1'h0;
      write_enable_data_log_force[4473] <= 1'h0;
      write_enable_data_log_force[4474] <= 1'h0;
      write_enable_data_log_force[4475] <= 1'h0;
      write_enable_data_log_force[4476] <= 1'h0;
      write_enable_data_log_force[4477] <= 1'h0;
      write_enable_data_log_force[4478] <= 1'h0;
      write_enable_data_log_force[4479] <= 1'h0;
      write_enable_data_log_force[4480] <= 1'h0;
      write_enable_data_log_force[4481] <= 1'h0;
      write_enable_data_log_force[4482] <= 1'h0;
      write_enable_data_log_force[4483] <= 1'h0;
      write_enable_data_log_force[4484] <= 1'h0;
      write_enable_data_log_force[4485] <= 1'h0;
      write_enable_data_log_force[4486] <= 1'h0;
      write_enable_data_log_force[4487] <= 1'h0;
      write_enable_data_log_force[4488] <= 1'h0;
      write_enable_data_log_force[4489] <= 1'h0;
      write_enable_data_log_force[4490] <= 1'h0;
      write_enable_data_log_force[4491] <= 1'h0;
      write_enable_data_log_force[4492] <= 1'h0;
      write_enable_data_log_force[4493] <= 1'h0;
      write_enable_data_log_force[4494] <= 1'h0;
      write_enable_data_log_force[4495] <= 1'h0;
      write_enable_data_log_force[4496] <= 1'h0;
      write_enable_data_log_force[4497] <= 1'h0;
      write_enable_data_log_force[4498] <= 1'h0;
      write_enable_data_log_force[4499] <= 1'h0;
      write_enable_data_log_force[4500] <= 1'h0;
      write_enable_data_log_force[4501] <= 1'h0;
      write_enable_data_log_force[4502] <= 1'h0;
      write_enable_data_log_force[4503] <= 1'h0;
      write_enable_data_log_force[4504] <= 1'h0;
      write_enable_data_log_force[4505] <= 1'h0;
      write_enable_data_log_force[4506] <= 1'h0;
      write_enable_data_log_force[4507] <= 1'h0;
      write_enable_data_log_force[4508] <= 1'h0;
      write_enable_data_log_force[4509] <= 1'h0;
      write_enable_data_log_force[4510] <= 1'h0;
      write_enable_data_log_force[4511] <= 1'h0;
      write_enable_data_log_force[4512] <= 1'h0;
      write_enable_data_log_force[4513] <= 1'h0;
      write_enable_data_log_force[4514] <= 1'h0;
      write_enable_data_log_force[4515] <= 1'h0;
      write_enable_data_log_force[4516] <= 1'h0;
      write_enable_data_log_force[4517] <= 1'h0;
      write_enable_data_log_force[4518] <= 1'h0;
      write_enable_data_log_force[4519] <= 1'h0;
      write_enable_data_log_force[4520] <= 1'h0;
      write_enable_data_log_force[4521] <= 1'h0;
      write_enable_data_log_force[4522] <= 1'h0;
      write_enable_data_log_force[4523] <= 1'h0;
      write_enable_data_log_force[4524] <= 1'h0;
      write_enable_data_log_force[4525] <= 1'h0;
      write_enable_data_log_force[4526] <= 1'h0;
      write_enable_data_log_force[4527] <= 1'h0;
      write_enable_data_log_force[4528] <= 1'h0;
      write_enable_data_log_force[4529] <= 1'h0;
      write_enable_data_log_force[4530] <= 1'h0;
      write_enable_data_log_force[4531] <= 1'h0;
      write_enable_data_log_force[4532] <= 1'h0;
      write_enable_data_log_force[4533] <= 1'h0;
      write_enable_data_log_force[4534] <= 1'h0;
      write_enable_data_log_force[4535] <= 1'h0;
      write_enable_data_log_force[4536] <= 1'h0;
      write_enable_data_log_force[4537] <= 1'h0;
      write_enable_data_log_force[4538] <= 1'h0;
      write_enable_data_log_force[4539] <= 1'h0;
      write_enable_data_log_force[4540] <= 1'h0;
      write_enable_data_log_force[4541] <= 1'h0;
      write_enable_data_log_force[4542] <= 1'h0;
      write_enable_data_log_force[4543] <= 1'h0;
      write_enable_data_log_force[4544] <= 1'h0;
      write_enable_data_log_force[4545] <= 1'h0;
      write_enable_data_log_force[4546] <= 1'h0;
      write_enable_data_log_force[4547] <= 1'h0;
      write_enable_data_log_force[4548] <= 1'h0;
      write_enable_data_log_force[4549] <= 1'h0;
      write_enable_data_log_force[4550] <= 1'h0;
      write_enable_data_log_force[4551] <= 1'h0;
      write_enable_data_log_force[4552] <= 1'h0;
      write_enable_data_log_force[4553] <= 1'h0;
      write_enable_data_log_force[4554] <= 1'h0;
      write_enable_data_log_force[4555] <= 1'h0;
      write_enable_data_log_force[4556] <= 1'h0;
      write_enable_data_log_force[4557] <= 1'h0;
      write_enable_data_log_force[4558] <= 1'h0;
      write_enable_data_log_force[4559] <= 1'h0;
      write_enable_data_log_force[4560] <= 1'h0;
      write_enable_data_log_force[4561] <= 1'h0;
      write_enable_data_log_force[4562] <= 1'h0;
      write_enable_data_log_force[4563] <= 1'h0;
      write_enable_data_log_force[4564] <= 1'h0;
      write_enable_data_log_force[4565] <= 1'h0;
      write_enable_data_log_force[4566] <= 1'h0;
      write_enable_data_log_force[4567] <= 1'h0;
      write_enable_data_log_force[4568] <= 1'h0;
      write_enable_data_log_force[4569] <= 1'h0;
      write_enable_data_log_force[4570] <= 1'h0;
      write_enable_data_log_force[4571] <= 1'h0;
      write_enable_data_log_force[4572] <= 1'h0;
      write_enable_data_log_force[4573] <= 1'h0;
      write_enable_data_log_force[4574] <= 1'h0;
      write_enable_data_log_force[4575] <= 1'h0;
      write_enable_data_log_force[4576] <= 1'h0;
      write_enable_data_log_force[4577] <= 1'h0;
      write_enable_data_log_force[4578] <= 1'h0;
      write_enable_data_log_force[4579] <= 1'h0;
      write_enable_data_log_force[4580] <= 1'h0;
      write_enable_data_log_force[4581] <= 1'h0;
      write_enable_data_log_force[4582] <= 1'h0;
      write_enable_data_log_force[4583] <= 1'h0;
      write_enable_data_log_force[4584] <= 1'h0;
      write_enable_data_log_force[4585] <= 1'h0;
      write_enable_data_log_force[4586] <= 1'h0;
      write_enable_data_log_force[4587] <= 1'h0;
      write_enable_data_log_force[4588] <= 1'h0;
      write_enable_data_log_force[4589] <= 1'h0;
      write_enable_data_log_force[4590] <= 1'h0;
      write_enable_data_log_force[4591] <= 1'h0;
      write_enable_data_log_force[4592] <= 1'h0;
      write_enable_data_log_force[4593] <= 1'h0;
      write_enable_data_log_force[4594] <= 1'h0;
      write_enable_data_log_force[4595] <= 1'h0;
      write_enable_data_log_force[4596] <= 1'h0;
      write_enable_data_log_force[4597] <= 1'h0;
      write_enable_data_log_force[4598] <= 1'h0;
      write_enable_data_log_force[4599] <= 1'h0;
      write_enable_data_log_force[4600] <= 1'h0;
      write_enable_data_log_force[4601] <= 1'h0;
      write_enable_data_log_force[4602] <= 1'h0;
      write_enable_data_log_force[4603] <= 1'h0;
      write_enable_data_log_force[4604] <= 1'h0;
      write_enable_data_log_force[4605] <= 1'h0;
      write_enable_data_log_force[4606] <= 1'h0;
      write_enable_data_log_force[4607] <= 1'h0;
      write_enable_data_log_force[4608] <= 1'h0;
      write_enable_data_log_force[4609] <= 1'h0;
      write_enable_data_log_force[4610] <= 1'h0;
      write_enable_data_log_force[4611] <= 1'h0;
      write_enable_data_log_force[4612] <= 1'h0;
      write_enable_data_log_force[4613] <= 1'h0;
      write_enable_data_log_force[4614] <= 1'h0;
      write_enable_data_log_force[4615] <= 1'h0;
      write_enable_data_log_force[4616] <= 1'h0;
      write_enable_data_log_force[4617] <= 1'h0;
      write_enable_data_log_force[4618] <= 1'h0;
      write_enable_data_log_force[4619] <= 1'h0;
      write_enable_data_log_force[4620] <= 1'h0;
      write_enable_data_log_force[4621] <= 1'h0;
      write_enable_data_log_force[4622] <= 1'h0;
      write_enable_data_log_force[4623] <= 1'h0;
      write_enable_data_log_force[4624] <= 1'h0;
      write_enable_data_log_force[4625] <= 1'h0;
      write_enable_data_log_force[4626] <= 1'h0;
      write_enable_data_log_force[4627] <= 1'h0;
      write_enable_data_log_force[4628] <= 1'h0;
      write_enable_data_log_force[4629] <= 1'h0;
      write_enable_data_log_force[4630] <= 1'h0;
      write_enable_data_log_force[4631] <= 1'h0;
      write_enable_data_log_force[4632] <= 1'h0;
      write_enable_data_log_force[4633] <= 1'h0;
      write_enable_data_log_force[4634] <= 1'h0;
      write_enable_data_log_force[4635] <= 1'h0;
      write_enable_data_log_force[4636] <= 1'h0;
      write_enable_data_log_force[4637] <= 1'h0;
      write_enable_data_log_force[4638] <= 1'h0;
      write_enable_data_log_force[4639] <= 1'h0;
      write_enable_data_log_force[4640] <= 1'h0;
      write_enable_data_log_force[4641] <= 1'h0;
      write_enable_data_log_force[4642] <= 1'h0;
      write_enable_data_log_force[4643] <= 1'h0;
      write_enable_data_log_force[4644] <= 1'h0;
      write_enable_data_log_force[4645] <= 1'h0;
      write_enable_data_log_force[4646] <= 1'h0;
      write_enable_data_log_force[4647] <= 1'h0;
      write_enable_data_log_force[4648] <= 1'h0;
      write_enable_data_log_force[4649] <= 1'h0;
      write_enable_data_log_force[4650] <= 1'h0;
      write_enable_data_log_force[4651] <= 1'h0;
      write_enable_data_log_force[4652] <= 1'h0;
      write_enable_data_log_force[4653] <= 1'h0;
      write_enable_data_log_force[4654] <= 1'h0;
      write_enable_data_log_force[4655] <= 1'h0;
      write_enable_data_log_force[4656] <= 1'h0;
      write_enable_data_log_force[4657] <= 1'h0;
      write_enable_data_log_force[4658] <= 1'h0;
      write_enable_data_log_force[4659] <= 1'h0;
      write_enable_data_log_force[4660] <= 1'h0;
      write_enable_data_log_force[4661] <= 1'h0;
      write_enable_data_log_force[4662] <= 1'h0;
      write_enable_data_log_force[4663] <= 1'h0;
      write_enable_data_log_force[4664] <= 1'h0;
      write_enable_data_log_force[4665] <= 1'h0;
      write_enable_data_log_force[4666] <= 1'h0;
      write_enable_data_log_force[4667] <= 1'h0;
      write_enable_data_log_force[4668] <= 1'h0;
      write_enable_data_log_force[4669] <= 1'h0;
      write_enable_data_log_force[4670] <= 1'h0;
      write_enable_data_log_force[4671] <= 1'h0;
      write_enable_data_log_force[4672] <= 1'h0;
      write_enable_data_log_force[4673] <= 1'h0;
      write_enable_data_log_force[4674] <= 1'h0;
      write_enable_data_log_force[4675] <= 1'h0;
      write_enable_data_log_force[4676] <= 1'h0;
      write_enable_data_log_force[4677] <= 1'h0;
      write_enable_data_log_force[4678] <= 1'h0;
      write_enable_data_log_force[4679] <= 1'h0;
      write_enable_data_log_force[4680] <= 1'h0;
      write_enable_data_log_force[4681] <= 1'h0;
      write_enable_data_log_force[4682] <= 1'h0;
      write_enable_data_log_force[4683] <= 1'h0;
      write_enable_data_log_force[4684] <= 1'h0;
      write_enable_data_log_force[4685] <= 1'h0;
      write_enable_data_log_force[4686] <= 1'h0;
      write_enable_data_log_force[4687] <= 1'h0;
      write_enable_data_log_force[4688] <= 1'h0;
      write_enable_data_log_force[4689] <= 1'h0;
      write_enable_data_log_force[4690] <= 1'h0;
      write_enable_data_log_force[4691] <= 1'h0;
      write_enable_data_log_force[4692] <= 1'h0;
      write_enable_data_log_force[4693] <= 1'h0;
      write_enable_data_log_force[4694] <= 1'h0;
      write_enable_data_log_force[4695] <= 1'h0;
      write_enable_data_log_force[4696] <= 1'h0;
      write_enable_data_log_force[4697] <= 1'h0;
      write_enable_data_log_force[4698] <= 1'h0;
      write_enable_data_log_force[4699] <= 1'h0;
      write_enable_data_log_force[4700] <= 1'h0;
      write_enable_data_log_force[4701] <= 1'h0;
      write_enable_data_log_force[4702] <= 1'h0;
      write_enable_data_log_force[4703] <= 1'h0;
      write_enable_data_log_force[4704] <= 1'h0;
      write_enable_data_log_force[4705] <= 1'h0;
      write_enable_data_log_force[4706] <= 1'h0;
      write_enable_data_log_force[4707] <= 1'h0;
      write_enable_data_log_force[4708] <= 1'h0;
      write_enable_data_log_force[4709] <= 1'h0;
      write_enable_data_log_force[4710] <= 1'h0;
      write_enable_data_log_force[4711] <= 1'h0;
      write_enable_data_log_force[4712] <= 1'h0;
      write_enable_data_log_force[4713] <= 1'h0;
      write_enable_data_log_force[4714] <= 1'h0;
      write_enable_data_log_force[4715] <= 1'h0;
      write_enable_data_log_force[4716] <= 1'h0;
      write_enable_data_log_force[4717] <= 1'h0;
      write_enable_data_log_force[4718] <= 1'h0;
      write_enable_data_log_force[4719] <= 1'h0;
      write_enable_data_log_force[4720] <= 1'h0;
      write_enable_data_log_force[4721] <= 1'h0;
      write_enable_data_log_force[4722] <= 1'h0;
      write_enable_data_log_force[4723] <= 1'h0;
      write_enable_data_log_force[4724] <= 1'h0;
      write_enable_data_log_force[4725] <= 1'h0;
      write_enable_data_log_force[4726] <= 1'h0;
      write_enable_data_log_force[4727] <= 1'h0;
      write_enable_data_log_force[4728] <= 1'h0;
      write_enable_data_log_force[4729] <= 1'h0;
      write_enable_data_log_force[4730] <= 1'h0;
      write_enable_data_log_force[4731] <= 1'h0;
      write_enable_data_log_force[4732] <= 1'h0;
      write_enable_data_log_force[4733] <= 1'h0;
      write_enable_data_log_force[4734] <= 1'h0;
      write_enable_data_log_force[4735] <= 1'h0;
      write_enable_data_log_force[4736] <= 1'h0;
      write_enable_data_log_force[4737] <= 1'h0;
      write_enable_data_log_force[4738] <= 1'h0;
      write_enable_data_log_force[4739] <= 1'h0;
      write_enable_data_log_force[4740] <= 1'h0;
      write_enable_data_log_force[4741] <= 1'h0;
      write_enable_data_log_force[4742] <= 1'h0;
      write_enable_data_log_force[4743] <= 1'h0;
      write_enable_data_log_force[4744] <= 1'h0;
      write_enable_data_log_force[4745] <= 1'h0;
      write_enable_data_log_force[4746] <= 1'h0;
      write_enable_data_log_force[4747] <= 1'h0;
      write_enable_data_log_force[4748] <= 1'h0;
      write_enable_data_log_force[4749] <= 1'h0;
      write_enable_data_log_force[4750] <= 1'h0;
      write_enable_data_log_force[4751] <= 1'h0;
      write_enable_data_log_force[4752] <= 1'h0;
      write_enable_data_log_force[4753] <= 1'h0;
      write_enable_data_log_force[4754] <= 1'h0;
      write_enable_data_log_force[4755] <= 1'h0;
      write_enable_data_log_force[4756] <= 1'h0;
      write_enable_data_log_force[4757] <= 1'h0;
      write_enable_data_log_force[4758] <= 1'h0;
      write_enable_data_log_force[4759] <= 1'h0;
      write_enable_data_log_force[4760] <= 1'h0;
      write_enable_data_log_force[4761] <= 1'h0;
      write_enable_data_log_force[4762] <= 1'h0;
      write_enable_data_log_force[4763] <= 1'h0;
      write_enable_data_log_force[4764] <= 1'h0;
      write_enable_data_log_force[4765] <= 1'h0;
      write_enable_data_log_force[4766] <= 1'h0;
      write_enable_data_log_force[4767] <= 1'h0;
      write_enable_data_log_force[4768] <= 1'h0;
      write_enable_data_log_force[4769] <= 1'h0;
      write_enable_data_log_force[4770] <= 1'h0;
      write_enable_data_log_force[4771] <= 1'h0;
      write_enable_data_log_force[4772] <= 1'h0;
      write_enable_data_log_force[4773] <= 1'h0;
      write_enable_data_log_force[4774] <= 1'h0;
      write_enable_data_log_force[4775] <= 1'h0;
      write_enable_data_log_force[4776] <= 1'h0;
      write_enable_data_log_force[4777] <= 1'h0;
      write_enable_data_log_force[4778] <= 1'h0;
      write_enable_data_log_force[4779] <= 1'h0;
      write_enable_data_log_force[4780] <= 1'h0;
      write_enable_data_log_force[4781] <= 1'h0;
      write_enable_data_log_force[4782] <= 1'h0;
      write_enable_data_log_force[4783] <= 1'h0;
      write_enable_data_log_force[4784] <= 1'h0;
      write_enable_data_log_force[4785] <= 1'h0;
      write_enable_data_log_force[4786] <= 1'h0;
      write_enable_data_log_force[4787] <= 1'h0;
      write_enable_data_log_force[4788] <= 1'h0;
      write_enable_data_log_force[4789] <= 1'h0;
      write_enable_data_log_force[4790] <= 1'h0;
      write_enable_data_log_force[4791] <= 1'h0;
      write_enable_data_log_force[4792] <= 1'h0;
      write_enable_data_log_force[4793] <= 1'h0;
      write_enable_data_log_force[4794] <= 1'h0;
      write_enable_data_log_force[4795] <= 1'h0;
      write_enable_data_log_force[4796] <= 1'h0;
      write_enable_data_log_force[4797] <= 1'h0;
      write_enable_data_log_force[4798] <= 1'h0;
      write_enable_data_log_force[4799] <= 1'h0;
      write_enable_data_log_force[4800] <= 1'h0;
      write_enable_data_log_force[4801] <= 1'h0;
      write_enable_data_log_force[4802] <= 1'h0;
      write_enable_data_log_force[4803] <= 1'h0;
      write_enable_data_log_force[4804] <= 1'h0;
      write_enable_data_log_force[4805] <= 1'h0;
      write_enable_data_log_force[4806] <= 1'h0;
      write_enable_data_log_force[4807] <= 1'h0;
      write_enable_data_log_force[4808] <= 1'h0;
      write_enable_data_log_force[4809] <= 1'h0;
      write_enable_data_log_force[4810] <= 1'h0;
      write_enable_data_log_force[4811] <= 1'h0;
      write_enable_data_log_force[4812] <= 1'h0;
      write_enable_data_log_force[4813] <= 1'h0;
      write_enable_data_log_force[4814] <= 1'h0;
      write_enable_data_log_force[4815] <= 1'h0;
      write_enable_data_log_force[4816] <= 1'h0;
      write_enable_data_log_force[4817] <= 1'h0;
      write_enable_data_log_force[4818] <= 1'h0;
      write_enable_data_log_force[4819] <= 1'h0;
      write_enable_data_log_force[4820] <= 1'h0;
      write_enable_data_log_force[4821] <= 1'h0;
      write_enable_data_log_force[4822] <= 1'h0;
      write_enable_data_log_force[4823] <= 1'h0;
      write_enable_data_log_force[4824] <= 1'h0;
      write_enable_data_log_force[4825] <= 1'h0;
      write_enable_data_log_force[4826] <= 1'h0;
      write_enable_data_log_force[4827] <= 1'h0;
      write_enable_data_log_force[4828] <= 1'h0;
      write_enable_data_log_force[4829] <= 1'h0;
      write_enable_data_log_force[4830] <= 1'h0;
      write_enable_data_log_force[4831] <= 1'h0;
      write_enable_data_log_force[4832] <= 1'h0;
      write_enable_data_log_force[4833] <= 1'h0;
      write_enable_data_log_force[4834] <= 1'h0;
      write_enable_data_log_force[4835] <= 1'h0;
      write_enable_data_log_force[4836] <= 1'h0;
      write_enable_data_log_force[4837] <= 1'h0;
      write_enable_data_log_force[4838] <= 1'h0;
      write_enable_data_log_force[4839] <= 1'h0;
      write_enable_data_log_force[4840] <= 1'h0;
      write_enable_data_log_force[4841] <= 1'h0;
      write_enable_data_log_force[4842] <= 1'h0;
      write_enable_data_log_force[4843] <= 1'h0;
      write_enable_data_log_force[4844] <= 1'h0;
      write_enable_data_log_force[4845] <= 1'h0;
      write_enable_data_log_force[4846] <= 1'h0;
      write_enable_data_log_force[4847] <= 1'h0;
      write_enable_data_log_force[4848] <= 1'h0;
      write_enable_data_log_force[4849] <= 1'h0;
      write_enable_data_log_force[4850] <= 1'h0;
      write_enable_data_log_force[4851] <= 1'h0;
      write_enable_data_log_force[4852] <= 1'h0;
      write_enable_data_log_force[4853] <= 1'h0;
      write_enable_data_log_force[4854] <= 1'h0;
      write_enable_data_log_force[4855] <= 1'h0;
      write_enable_data_log_force[4856] <= 1'h0;
      write_enable_data_log_force[4857] <= 1'h0;
      write_enable_data_log_force[4858] <= 1'h0;
      write_enable_data_log_force[4859] <= 1'h0;
      write_enable_data_log_force[4860] <= 1'h0;
      write_enable_data_log_force[4861] <= 1'h0;
      write_enable_data_log_force[4862] <= 1'h0;
      write_enable_data_log_force[4863] <= 1'h0;
      write_enable_data_log_force[4864] <= 1'h0;
      write_enable_data_log_force[4865] <= 1'h0;
      write_enable_data_log_force[4866] <= 1'h0;
      write_enable_data_log_force[4867] <= 1'h0;
      write_enable_data_log_force[4868] <= 1'h0;
      write_enable_data_log_force[4869] <= 1'h0;
      write_enable_data_log_force[4870] <= 1'h0;
      write_enable_data_log_force[4871] <= 1'h0;
      write_enable_data_log_force[4872] <= 1'h0;
      write_enable_data_log_force[4873] <= 1'h0;
      write_enable_data_log_force[4874] <= 1'h0;
      write_enable_data_log_force[4875] <= 1'h0;
      write_enable_data_log_force[4876] <= 1'h0;
      write_enable_data_log_force[4877] <= 1'h0;
      write_enable_data_log_force[4878] <= 1'h0;
      write_enable_data_log_force[4879] <= 1'h0;
      write_enable_data_log_force[4880] <= 1'h0;
      write_enable_data_log_force[4881] <= 1'h0;
      write_enable_data_log_force[4882] <= 1'h0;
      write_enable_data_log_force[4883] <= 1'h0;
      write_enable_data_log_force[4884] <= 1'h0;
      write_enable_data_log_force[4885] <= 1'h0;
      write_enable_data_log_force[4886] <= 1'h0;
      write_enable_data_log_force[4887] <= 1'h0;
      write_enable_data_log_force[4888] <= 1'h0;
      write_enable_data_log_force[4889] <= 1'h0;
      write_enable_data_log_force[4890] <= 1'h0;
      write_enable_data_log_force[4891] <= 1'h0;
      write_enable_data_log_force[4892] <= 1'h0;
      write_enable_data_log_force[4893] <= 1'h0;
      write_enable_data_log_force[4894] <= 1'h0;
      write_enable_data_log_force[4895] <= 1'h0;
      write_enable_data_log_force[4896] <= 1'h0;
      write_enable_data_log_force[4897] <= 1'h0;
      write_enable_data_log_force[4898] <= 1'h0;
      write_enable_data_log_force[4899] <= 1'h0;
      write_enable_data_log_force[4900] <= 1'h0;
      write_enable_data_log_force[4901] <= 1'h0;
      write_enable_data_log_force[4902] <= 1'h0;
      write_enable_data_log_force[4903] <= 1'h0;
      write_enable_data_log_force[4904] <= 1'h0;
      write_enable_data_log_force[4905] <= 1'h0;
      write_enable_data_log_force[4906] <= 1'h0;
      write_enable_data_log_force[4907] <= 1'h0;
      write_enable_data_log_force[4908] <= 1'h0;
      write_enable_data_log_force[4909] <= 1'h0;
      write_enable_data_log_force[4910] <= 1'h0;
      write_enable_data_log_force[4911] <= 1'h0;
      write_enable_data_log_force[4912] <= 1'h0;
      write_enable_data_log_force[4913] <= 1'h0;
      write_enable_data_log_force[4914] <= 1'h0;
      write_enable_data_log_force[4915] <= 1'h0;
      write_enable_data_log_force[4916] <= 1'h0;
      write_enable_data_log_force[4917] <= 1'h0;
      write_enable_data_log_force[4918] <= 1'h0;
      write_enable_data_log_force[4919] <= 1'h0;
      write_enable_data_log_force[4920] <= 1'h0;
      write_enable_data_log_force[4921] <= 1'h0;
      write_enable_data_log_force[4922] <= 1'h0;
      write_enable_data_log_force[4923] <= 1'h0;
      write_enable_data_log_force[4924] <= 1'h0;
      write_enable_data_log_force[4925] <= 1'h0;
      write_enable_data_log_force[4926] <= 1'h0;
      write_enable_data_log_force[4927] <= 1'h0;
      write_enable_data_log_force[4928] <= 1'h0;
      write_enable_data_log_force[4929] <= 1'h0;
      write_enable_data_log_force[4930] <= 1'h0;
      write_enable_data_log_force[4931] <= 1'h0;
      write_enable_data_log_force[4932] <= 1'h0;
      write_enable_data_log_force[4933] <= 1'h0;
      write_enable_data_log_force[4934] <= 1'h0;
      write_enable_data_log_force[4935] <= 1'h0;
      write_enable_data_log_force[4936] <= 1'h0;
      write_enable_data_log_force[4937] <= 1'h0;
      write_enable_data_log_force[4938] <= 1'h0;
      write_enable_data_log_force[4939] <= 1'h0;
      write_enable_data_log_force[4940] <= 1'h0;
      write_enable_data_log_force[4941] <= 1'h0;
      write_enable_data_log_force[4942] <= 1'h0;
      write_enable_data_log_force[4943] <= 1'h0;
      write_enable_data_log_force[4944] <= 1'h0;
      write_enable_data_log_force[4945] <= 1'h0;
      write_enable_data_log_force[4946] <= 1'h0;
      write_enable_data_log_force[4947] <= 1'h0;
      write_enable_data_log_force[4948] <= 1'h0;
      write_enable_data_log_force[4949] <= 1'h0;
      write_enable_data_log_force[4950] <= 1'h0;
      write_enable_data_log_force[4951] <= 1'h0;
      write_enable_data_log_force[4952] <= 1'h0;
      write_enable_data_log_force[4953] <= 1'h0;
      write_enable_data_log_force[4954] <= 1'h0;
      write_enable_data_log_force[4955] <= 1'h0;
      write_enable_data_log_force[4956] <= 1'h0;
      write_enable_data_log_force[4957] <= 1'h0;
      write_enable_data_log_force[4958] <= 1'h0;
      write_enable_data_log_force[4959] <= 1'h0;
      write_enable_data_log_force[4960] <= 1'h0;
      write_enable_data_log_force[4961] <= 1'h0;
      write_enable_data_log_force[4962] <= 1'h0;
      write_enable_data_log_force[4963] <= 1'h0;
      write_enable_data_log_force[4964] <= 1'h0;
      write_enable_data_log_force[4965] <= 1'h0;
      write_enable_data_log_force[4966] <= 1'h0;
      write_enable_data_log_force[4967] <= 1'h0;
      write_enable_data_log_force[4968] <= 1'h0;
      write_enable_data_log_force[4969] <= 1'h0;
      write_enable_data_log_force[4970] <= 1'h0;
      write_enable_data_log_force[4971] <= 1'h0;
      write_enable_data_log_force[4972] <= 1'h0;
      write_enable_data_log_force[4973] <= 1'h0;
      write_enable_data_log_force[4974] <= 1'h0;
      write_enable_data_log_force[4975] <= 1'h0;
      write_enable_data_log_force[4976] <= 1'h0;
      write_enable_data_log_force[4977] <= 1'h0;
      write_enable_data_log_force[4978] <= 1'h0;
      write_enable_data_log_force[4979] <= 1'h0;
      write_enable_data_log_force[4980] <= 1'h0;
      write_enable_data_log_force[4981] <= 1'h0;
      write_enable_data_log_force[4982] <= 1'h0;
      write_enable_data_log_force[4983] <= 1'h0;
      write_enable_data_log_force[4984] <= 1'h0;
      write_enable_data_log_force[4985] <= 1'h0;
      write_enable_data_log_force[4986] <= 1'h0;
      write_enable_data_log_force[4987] <= 1'h0;
      write_enable_data_log_force[4988] <= 1'h0;
      write_enable_data_log_force[4989] <= 1'h0;
      write_enable_data_log_force[4990] <= 1'h0;
      write_enable_data_log_force[4991] <= 1'h0;
      write_enable_data_log_force[4992] <= 1'h0;
      write_enable_data_log_force[4993] <= 1'h0;
      write_enable_data_log_force[4994] <= 1'h0;
      write_enable_data_log_force[4995] <= 1'h0;
      write_enable_data_log_force[4996] <= 1'h0;
      write_enable_data_log_force[4997] <= 1'h0;
      write_enable_data_log_force[4998] <= 1'h0;
      write_enable_data_log_force[4999] <= 1'h0;
      write_enable_data_log_force[5000] <= 1'h0;
      write_enable_data_log_force[5001] <= 1'h0;
      write_enable_data_log_force[5002] <= 1'h0;
      write_enable_data_log_force[5003] <= 1'h0;
      write_enable_data_log_force[5004] <= 1'h0;
      write_enable_data_log_force[5005] <= 1'h0;
      write_enable_data_log_force[5006] <= 1'h0;
      write_enable_data_log_force[5007] <= 1'h0;
      write_enable_data_log_force[5008] <= 1'h0;
      write_enable_data_log_force[5009] <= 1'h0;
      write_enable_data_log_force[5010] <= 1'h0;
      write_enable_data_log_force[5011] <= 1'h0;
      write_enable_data_log_force[5012] <= 1'h0;
      write_enable_data_log_force[5013] <= 1'h0;
      write_enable_data_log_force[5014] <= 1'h0;
      write_enable_data_log_force[5015] <= 1'h0;
      write_enable_data_log_force[5016] <= 1'h0;
      write_enable_data_log_force[5017] <= 1'h0;
      write_enable_data_log_force[5018] <= 1'h0;
      write_enable_data_log_force[5019] <= 1'h0;
      write_enable_data_log_force[5020] <= 1'h0;
      write_enable_data_log_force[5021] <= 1'h0;
      write_enable_data_log_force[5022] <= 1'h0;
      write_enable_data_log_force[5023] <= 1'h0;
      write_enable_data_log_force[5024] <= 1'h0;
      write_enable_data_log_force[5025] <= 1'h0;
      write_enable_data_log_force[5026] <= 1'h0;
      write_enable_data_log_force[5027] <= 1'h0;
      write_enable_data_log_force[5028] <= 1'h0;
      write_enable_data_log_force[5029] <= 1'h0;
      write_enable_data_log_force[5030] <= 1'h0;
      write_enable_data_log_force[5031] <= 1'h0;
      write_enable_data_log_force[5032] <= 1'h0;
      write_enable_data_log_force[5033] <= 1'h0;
      write_enable_data_log_force[5034] <= 1'h0;
      write_enable_data_log_force[5035] <= 1'h0;
      write_enable_data_log_force[5036] <= 1'h0;
      write_enable_data_log_force[5037] <= 1'h0;
      write_enable_data_log_force[5038] <= 1'h0;
      write_enable_data_log_force[5039] <= 1'h0;
      write_enable_data_log_force[5040] <= 1'h0;
      write_enable_data_log_force[5041] <= 1'h0;
      write_enable_data_log_force[5042] <= 1'h0;
      write_enable_data_log_force[5043] <= 1'h0;
      write_enable_data_log_force[5044] <= 1'h0;
      write_enable_data_log_force[5045] <= 1'h0;
      write_enable_data_log_force[5046] <= 1'h0;
      write_enable_data_log_force[5047] <= 1'h0;
      write_enable_data_log_force[5048] <= 1'h0;
      write_enable_data_log_force[5049] <= 1'h0;
      write_enable_data_log_force[5050] <= 1'h0;
      write_enable_data_log_force[5051] <= 1'h0;
      write_enable_data_log_force[5052] <= 1'h0;
      write_enable_data_log_force[5053] <= 1'h0;
      write_enable_data_log_force[5054] <= 1'h0;
      write_enable_data_log_force[5055] <= 1'h0;
      write_enable_data_log_force[5056] <= 1'h0;
      write_enable_data_log_force[5057] <= 1'h0;
      write_enable_data_log_force[5058] <= 1'h0;
      write_enable_data_log_force[5059] <= 1'h0;
      write_enable_data_log_force[5060] <= 1'h0;
      write_enable_data_log_force[5061] <= 1'h0;
      write_enable_data_log_force[5062] <= 1'h0;
      write_enable_data_log_force[5063] <= 1'h0;
      write_enable_data_log_force[5064] <= 1'h0;
      write_enable_data_log_force[5065] <= 1'h0;
      write_enable_data_log_force[5066] <= 1'h0;
      write_enable_data_log_force[5067] <= 1'h0;
      write_enable_data_log_force[5068] <= 1'h0;
      write_enable_data_log_force[5069] <= 1'h0;
      write_enable_data_log_force[5070] <= 1'h0;
      write_enable_data_log_force[5071] <= 1'h0;
      write_enable_data_log_force[5072] <= 1'h0;
      write_enable_data_log_force[5073] <= 1'h0;
      write_enable_data_log_force[5074] <= 1'h0;
      write_enable_data_log_force[5075] <= 1'h0;
      write_enable_data_log_force[5076] <= 1'h0;
      write_enable_data_log_force[5077] <= 1'h0;
      write_enable_data_log_force[5078] <= 1'h0;
      write_enable_data_log_force[5079] <= 1'h0;
      write_enable_data_log_force[5080] <= 1'h0;
      write_enable_data_log_force[5081] <= 1'h0;
      write_enable_data_log_force[5082] <= 1'h0;
      write_enable_data_log_force[5083] <= 1'h0;
      write_enable_data_log_force[5084] <= 1'h0;
      write_enable_data_log_force[5085] <= 1'h0;
      write_enable_data_log_force[5086] <= 1'h0;
      write_enable_data_log_force[5087] <= 1'h0;
      write_enable_data_log_force[5088] <= 1'h0;
      write_enable_data_log_force[5089] <= 1'h0;
      write_enable_data_log_force[5090] <= 1'h0;
      write_enable_data_log_force[5091] <= 1'h0;
      write_enable_data_log_force[5092] <= 1'h0;
      write_enable_data_log_force[5093] <= 1'h0;
      write_enable_data_log_force[5094] <= 1'h0;
      write_enable_data_log_force[5095] <= 1'h0;
      write_enable_data_log_force[5096] <= 1'h0;
      write_enable_data_log_force[5097] <= 1'h0;
      write_enable_data_log_force[5098] <= 1'h0;
      write_enable_data_log_force[5099] <= 1'h0;
      write_enable_data_log_force[5100] <= 1'h0;
      write_enable_data_log_force[5101] <= 1'h0;
      write_enable_data_log_force[5102] <= 1'h0;
      write_enable_data_log_force[5103] <= 1'h0;
      write_enable_data_log_force[5104] <= 1'h0;
      write_enable_data_log_force[5105] <= 1'h0;
      write_enable_data_log_force[5106] <= 1'h0;
      write_enable_data_log_force[5107] <= 1'h0;
      write_enable_data_log_force[5108] <= 1'h0;
      write_enable_data_log_force[5109] <= 1'h0;
      write_enable_data_log_force[5110] <= 1'h0;
      write_enable_data_log_force[5111] <= 1'h0;
      write_enable_data_log_force[5112] <= 1'h0;
      write_enable_data_log_force[5113] <= 1'h0;
      write_enable_data_log_force[5114] <= 1'h0;
      write_enable_data_log_force[5115] <= 1'h0;
      write_enable_data_log_force[5116] <= 1'h0;
      write_enable_data_log_force[5117] <= 1'h0;
      write_enable_data_log_force[5118] <= 1'h0;
      write_enable_data_log_force[5119] <= 1'h0;
      write_enable_data_log_force[5120] <= 1'h0;
      write_enable_data_log_force[5121] <= 1'h0;
      write_enable_data_log_force[5122] <= 1'h0;
      write_enable_data_log_force[5123] <= 1'h0;
      write_enable_data_log_force[5124] <= 1'h0;
      write_enable_data_log_force[5125] <= 1'h0;
      write_enable_data_log_force[5126] <= 1'h0;
      write_enable_data_log_force[5127] <= 1'h0;
      write_enable_data_log_force[5128] <= 1'h0;
      write_enable_data_log_force[5129] <= 1'h0;
      write_enable_data_log_force[5130] <= 1'h0;
      write_enable_data_log_force[5131] <= 1'h0;
      write_enable_data_log_force[5132] <= 1'h0;
      write_enable_data_log_force[5133] <= 1'h0;
      write_enable_data_log_force[5134] <= 1'h0;
      write_enable_data_log_force[5135] <= 1'h0;
      write_enable_data_log_force[5136] <= 1'h0;
      write_enable_data_log_force[5137] <= 1'h0;
      write_enable_data_log_force[5138] <= 1'h0;
      write_enable_data_log_force[5139] <= 1'h0;
      write_enable_data_log_force[5140] <= 1'h0;
      write_enable_data_log_force[5141] <= 1'h0;
      write_enable_data_log_force[5142] <= 1'h0;
      write_enable_data_log_force[5143] <= 1'h0;
      write_enable_data_log_force[5144] <= 1'h0;
      write_enable_data_log_force[5145] <= 1'h0;
      write_enable_data_log_force[5146] <= 1'h0;
      write_enable_data_log_force[5147] <= 1'h0;
      write_enable_data_log_force[5148] <= 1'h0;
      write_enable_data_log_force[5149] <= 1'h0;
      write_enable_data_log_force[5150] <= 1'h0;
      write_enable_data_log_force[5151] <= 1'h0;
      write_enable_data_log_force[5152] <= 1'h0;
      write_enable_data_log_force[5153] <= 1'h0;
      write_enable_data_log_force[5154] <= 1'h0;
      write_enable_data_log_force[5155] <= 1'h0;
      write_enable_data_log_force[5156] <= 1'h0;
      write_enable_data_log_force[5157] <= 1'h0;
      write_enable_data_log_force[5158] <= 1'h0;
      write_enable_data_log_force[5159] <= 1'h0;
      write_enable_data_log_force[5160] <= 1'h0;
      write_enable_data_log_force[5161] <= 1'h0;
      write_enable_data_log_force[5162] <= 1'h0;
      write_enable_data_log_force[5163] <= 1'h0;
      write_enable_data_log_force[5164] <= 1'h0;
      write_enable_data_log_force[5165] <= 1'h0;
      write_enable_data_log_force[5166] <= 1'h0;
      write_enable_data_log_force[5167] <= 1'h0;
      write_enable_data_log_force[5168] <= 1'h0;
      write_enable_data_log_force[5169] <= 1'h0;
      write_enable_data_log_force[5170] <= 1'h0;
      write_enable_data_log_force[5171] <= 1'h0;
      write_enable_data_log_force[5172] <= 1'h0;
      write_enable_data_log_force[5173] <= 1'h0;
      write_enable_data_log_force[5174] <= 1'h0;
      write_enable_data_log_force[5175] <= 1'h0;
      write_enable_data_log_force[5176] <= 1'h0;
      write_enable_data_log_force[5177] <= 1'h0;
      write_enable_data_log_force[5178] <= 1'h0;
      write_enable_data_log_force[5179] <= 1'h0;
      write_enable_data_log_force[5180] <= 1'h0;
      write_enable_data_log_force[5181] <= 1'h0;
      write_enable_data_log_force[5182] <= 1'h0;
      write_enable_data_log_force[5183] <= 1'h0;
      write_enable_data_log_force[5184] <= 1'h0;
      write_enable_data_log_force[5185] <= 1'h0;
      write_enable_data_log_force[5186] <= 1'h0;
      write_enable_data_log_force[5187] <= 1'h0;
      write_enable_data_log_force[5188] <= 1'h0;
      write_enable_data_log_force[5189] <= 1'h0;
      write_enable_data_log_force[5190] <= 1'h0;
      write_enable_data_log_force[5191] <= 1'h0;
      write_enable_data_log_force[5192] <= 1'h0;
      write_enable_data_log_force[5193] <= 1'h0;
      write_enable_data_log_force[5194] <= 1'h0;
      write_enable_data_log_force[5195] <= 1'h0;
      write_enable_data_log_force[5196] <= 1'h0;
      write_enable_data_log_force[5197] <= 1'h0;
      write_enable_data_log_force[5198] <= 1'h0;
      write_enable_data_log_force[5199] <= 1'h0;
      write_enable_data_log_force[5200] <= 1'h0;
      write_enable_data_log_force[5201] <= 1'h0;
      write_enable_data_log_force[5202] <= 1'h0;
      write_enable_data_log_force[5203] <= 1'h0;
      write_enable_data_log_force[5204] <= 1'h0;
      write_enable_data_log_force[5205] <= 1'h0;
      write_enable_data_log_force[5206] <= 1'h0;
      write_enable_data_log_force[5207] <= 1'h0;
      write_enable_data_log_force[5208] <= 1'h0;
      write_enable_data_log_force[5209] <= 1'h0;
      write_enable_data_log_force[5210] <= 1'h0;
      write_enable_data_log_force[5211] <= 1'h0;
      write_enable_data_log_force[5212] <= 1'h0;
      write_enable_data_log_force[5213] <= 1'h0;
      write_enable_data_log_force[5214] <= 1'h0;
      write_enable_data_log_force[5215] <= 1'h0;
      write_enable_data_log_force[5216] <= 1'h0;
      write_enable_data_log_force[5217] <= 1'h0;
      write_enable_data_log_force[5218] <= 1'h0;
      write_enable_data_log_force[5219] <= 1'h0;
      write_enable_data_log_force[5220] <= 1'h0;
      write_enable_data_log_force[5221] <= 1'h0;
      write_enable_data_log_force[5222] <= 1'h0;
      write_enable_data_log_force[5223] <= 1'h0;
      write_enable_data_log_force[5224] <= 1'h0;
      write_enable_data_log_force[5225] <= 1'h0;
      write_enable_data_log_force[5226] <= 1'h0;
      write_enable_data_log_force[5227] <= 1'h0;
      write_enable_data_log_force[5228] <= 1'h0;
      write_enable_data_log_force[5229] <= 1'h0;
      write_enable_data_log_force[5230] <= 1'h0;
      write_enable_data_log_force[5231] <= 1'h0;
      write_enable_data_log_force[5232] <= 1'h0;
      write_enable_data_log_force[5233] <= 1'h0;
      write_enable_data_log_force[5234] <= 1'h0;
      write_enable_data_log_force[5235] <= 1'h0;
      write_enable_data_log_force[5236] <= 1'h0;
      write_enable_data_log_force[5237] <= 1'h0;
      write_enable_data_log_force[5238] <= 1'h0;
      write_enable_data_log_force[5239] <= 1'h0;
      write_enable_data_log_force[5240] <= 1'h0;
      write_enable_data_log_force[5241] <= 1'h0;
      write_enable_data_log_force[5242] <= 1'h0;
      write_enable_data_log_force[5243] <= 1'h0;
      write_enable_data_log_force[5244] <= 1'h0;
      write_enable_data_log_force[5245] <= 1'h0;
      write_enable_data_log_force[5246] <= 1'h0;
      write_enable_data_log_force[5247] <= 1'h0;
      write_enable_data_log_force[5248] <= 1'h0;
      write_enable_data_log_force[5249] <= 1'h0;
      write_enable_data_log_force[5250] <= 1'h0;
      write_enable_data_log_force[5251] <= 1'h0;
      write_enable_data_log_force[5252] <= 1'h0;
      write_enable_data_log_force[5253] <= 1'h0;
      write_enable_data_log_force[5254] <= 1'h0;
      write_enable_data_log_force[5255] <= 1'h0;
      write_enable_data_log_force[5256] <= 1'h0;
      write_enable_data_log_force[5257] <= 1'h0;
      write_enable_data_log_force[5258] <= 1'h0;
      write_enable_data_log_force[5259] <= 1'h0;
      write_enable_data_log_force[5260] <= 1'h0;
      write_enable_data_log_force[5261] <= 1'h0;
      write_enable_data_log_force[5262] <= 1'h0;
      write_enable_data_log_force[5263] <= 1'h0;
      write_enable_data_log_force[5264] <= 1'h0;
      write_enable_data_log_force[5265] <= 1'h0;
      write_enable_data_log_force[5266] <= 1'h0;
      write_enable_data_log_force[5267] <= 1'h0;
      write_enable_data_log_force[5268] <= 1'h0;
      write_enable_data_log_force[5269] <= 1'h0;
      write_enable_data_log_force[5270] <= 1'h0;
      write_enable_data_log_force[5271] <= 1'h0;
      write_enable_data_log_force[5272] <= 1'h0;
      write_enable_data_log_force[5273] <= 1'h0;
      write_enable_data_log_force[5274] <= 1'h0;
      write_enable_data_log_force[5275] <= 1'h0;
      write_enable_data_log_force[5276] <= 1'h0;
      write_enable_data_log_force[5277] <= 1'h0;
      write_enable_data_log_force[5278] <= 1'h0;
      write_enable_data_log_force[5279] <= 1'h0;
      write_enable_data_log_force[5280] <= 1'h0;
      write_enable_data_log_force[5281] <= 1'h0;
      write_enable_data_log_force[5282] <= 1'h0;
      write_enable_data_log_force[5283] <= 1'h0;
      write_enable_data_log_force[5284] <= 1'h0;
      write_enable_data_log_force[5285] <= 1'h0;
      write_enable_data_log_force[5286] <= 1'h0;
      write_enable_data_log_force[5287] <= 1'h0;
      write_enable_data_log_force[5288] <= 1'h0;
      write_enable_data_log_force[5289] <= 1'h0;
      write_enable_data_log_force[5290] <= 1'h0;
      write_enable_data_log_force[5291] <= 1'h0;
      write_enable_data_log_force[5292] <= 1'h0;
      write_enable_data_log_force[5293] <= 1'h0;
      write_enable_data_log_force[5294] <= 1'h0;
      write_enable_data_log_force[5295] <= 1'h0;
      write_enable_data_log_force[5296] <= 1'h0;
      write_enable_data_log_force[5297] <= 1'h0;
      write_enable_data_log_force[5298] <= 1'h0;
      write_enable_data_log_force[5299] <= 1'h0;
      write_enable_data_log_force[5300] <= 1'h0;
      write_enable_data_log_force[5301] <= 1'h0;
      write_enable_data_log_force[5302] <= 1'h0;
      write_enable_data_log_force[5303] <= 1'h0;
      write_enable_data_log_force[5304] <= 1'h0;
      write_enable_data_log_force[5305] <= 1'h0;
      write_enable_data_log_force[5306] <= 1'h0;
      write_enable_data_log_force[5307] <= 1'h0;
      write_enable_data_log_force[5308] <= 1'h0;
      write_enable_data_log_force[5309] <= 1'h0;
      write_enable_data_log_force[5310] <= 1'h0;
      write_enable_data_log_force[5311] <= 1'h0;
      write_enable_data_log_force[5312] <= 1'h0;
      write_enable_data_log_force[5313] <= 1'h0;
      write_enable_data_log_force[5314] <= 1'h0;
      write_enable_data_log_force[5315] <= 1'h0;
      write_enable_data_log_force[5316] <= 1'h0;
      write_enable_data_log_force[5317] <= 1'h0;
      write_enable_data_log_force[5318] <= 1'h0;
      write_enable_data_log_force[5319] <= 1'h0;
      write_enable_data_log_force[5320] <= 1'h0;
      write_enable_data_log_force[5321] <= 1'h0;
      write_enable_data_log_force[5322] <= 1'h0;
      write_enable_data_log_force[5323] <= 1'h0;
      write_enable_data_log_force[5324] <= 1'h0;
      write_enable_data_log_force[5325] <= 1'h0;
      write_enable_data_log_force[5326] <= 1'h0;
      write_enable_data_log_force[5327] <= 1'h0;
      write_enable_data_log_force[5328] <= 1'h0;
      write_enable_data_log_force[5329] <= 1'h0;
      write_enable_data_log_force[5330] <= 1'h0;
      write_enable_data_log_force[5331] <= 1'h0;
      write_enable_data_log_force[5332] <= 1'h0;
      write_enable_data_log_force[5333] <= 1'h0;
      write_enable_data_log_force[5334] <= 1'h0;
      write_enable_data_log_force[5335] <= 1'h0;
      write_enable_data_log_force[5336] <= 1'h0;
      write_enable_data_log_force[5337] <= 1'h0;
      write_enable_data_log_force[5338] <= 1'h0;
      write_enable_data_log_force[5339] <= 1'h0;
      write_enable_data_log_force[5340] <= 1'h0;
      write_enable_data_log_force[5341] <= 1'h0;
      write_enable_data_log_force[5342] <= 1'h0;
      write_enable_data_log_force[5343] <= 1'h0;
      write_enable_data_log_force[5344] <= 1'h0;
      write_enable_data_log_force[5345] <= 1'h0;
      write_enable_data_log_force[5346] <= 1'h0;
      write_enable_data_log_force[5347] <= 1'h0;
      write_enable_data_log_force[5348] <= 1'h0;
      write_enable_data_log_force[5349] <= 1'h0;
      write_enable_data_log_force[5350] <= 1'h0;
      write_enable_data_log_force[5351] <= 1'h0;
      write_enable_data_log_force[5352] <= 1'h0;
      write_enable_data_log_force[5353] <= 1'h0;
      write_enable_data_log_force[5354] <= 1'h0;
      write_enable_data_log_force[5355] <= 1'h0;
      write_enable_data_log_force[5356] <= 1'h0;
      write_enable_data_log_force[5357] <= 1'h0;
      write_enable_data_log_force[5358] <= 1'h0;
      write_enable_data_log_force[5359] <= 1'h0;
      write_enable_data_log_force[5360] <= 1'h0;
      write_enable_data_log_force[5361] <= 1'h0;
      write_enable_data_log_force[5362] <= 1'h0;
      write_enable_data_log_force[5363] <= 1'h0;
      write_enable_data_log_force[5364] <= 1'h0;
      write_enable_data_log_force[5365] <= 1'h0;
      write_enable_data_log_force[5366] <= 1'h0;
      write_enable_data_log_force[5367] <= 1'h0;
      write_enable_data_log_force[5368] <= 1'h0;
      write_enable_data_log_force[5369] <= 1'h0;
      write_enable_data_log_force[5370] <= 1'h0;
      write_enable_data_log_force[5371] <= 1'h0;
      write_enable_data_log_force[5372] <= 1'h0;
      write_enable_data_log_force[5373] <= 1'h0;
      write_enable_data_log_force[5374] <= 1'h0;
      write_enable_data_log_force[5375] <= 1'h0;
      write_enable_data_log_force[5376] <= 1'h0;
      write_enable_data_log_force[5377] <= 1'h0;
      write_enable_data_log_force[5378] <= 1'h0;
      write_enable_data_log_force[5379] <= 1'h0;
      write_enable_data_log_force[5380] <= 1'h0;
      write_enable_data_log_force[5381] <= 1'h0;
      write_enable_data_log_force[5382] <= 1'h0;
      write_enable_data_log_force[5383] <= 1'h0;
      write_enable_data_log_force[5384] <= 1'h0;
      write_enable_data_log_force[5385] <= 1'h0;
      write_enable_data_log_force[5386] <= 1'h0;
      write_enable_data_log_force[5387] <= 1'h0;
      write_enable_data_log_force[5388] <= 1'h0;
      write_enable_data_log_force[5389] <= 1'h0;
      write_enable_data_log_force[5390] <= 1'h0;
      write_enable_data_log_force[5391] <= 1'h0;
      write_enable_data_log_force[5392] <= 1'h0;
      write_enable_data_log_force[5393] <= 1'h0;
      write_enable_data_log_force[5394] <= 1'h0;
      write_enable_data_log_force[5395] <= 1'h0;
      write_enable_data_log_force[5396] <= 1'h0;
      write_enable_data_log_force[5397] <= 1'h0;
      write_enable_data_log_force[5398] <= 1'h0;
      write_enable_data_log_force[5399] <= 1'h0;
      write_enable_data_log_force[5400] <= 1'h0;
      write_enable_data_log_force[5401] <= 1'h0;
      write_enable_data_log_force[5402] <= 1'h0;
      write_enable_data_log_force[5403] <= 1'h0;
      write_enable_data_log_force[5404] <= 1'h0;
      write_enable_data_log_force[5405] <= 1'h0;
      write_enable_data_log_force[5406] <= 1'h0;
      write_enable_data_log_force[5407] <= 1'h0;
      write_enable_data_log_force[5408] <= 1'h0;
      write_enable_data_log_force[5409] <= 1'h0;
      write_enable_data_log_force[5410] <= 1'h0;
      write_enable_data_log_force[5411] <= 1'h0;
      write_enable_data_log_force[5412] <= 1'h0;
      write_enable_data_log_force[5413] <= 1'h0;
      write_enable_data_log_force[5414] <= 1'h0;
      write_enable_data_log_force[5415] <= 1'h0;
      write_enable_data_log_force[5416] <= 1'h0;
      write_enable_data_log_force[5417] <= 1'h0;
      write_enable_data_log_force[5418] <= 1'h0;
      write_enable_data_log_force[5419] <= 1'h0;
      write_enable_data_log_force[5420] <= 1'h0;
      write_enable_data_log_force[5421] <= 1'h0;
      write_enable_data_log_force[5422] <= 1'h0;
      write_enable_data_log_force[5423] <= 1'h0;
      write_enable_data_log_force[5424] <= 1'h0;
      write_enable_data_log_force[5425] <= 1'h0;
      write_enable_data_log_force[5426] <= 1'h0;
      write_enable_data_log_force[5427] <= 1'h0;
      write_enable_data_log_force[5428] <= 1'h0;
      write_enable_data_log_force[5429] <= 1'h0;
      write_enable_data_log_force[5430] <= 1'h0;
      write_enable_data_log_force[5431] <= 1'h0;
      write_enable_data_log_force[5432] <= 1'h0;
      write_enable_data_log_force[5433] <= 1'h0;
      write_enable_data_log_force[5434] <= 1'h0;
      write_enable_data_log_force[5435] <= 1'h0;
      write_enable_data_log_force[5436] <= 1'h0;
      write_enable_data_log_force[5437] <= 1'h0;
      write_enable_data_log_force[5438] <= 1'h0;
      write_enable_data_log_force[5439] <= 1'h0;
      write_enable_data_log_force[5440] <= 1'h0;
      write_enable_data_log_force[5441] <= 1'h0;
      write_enable_data_log_force[5442] <= 1'h0;
      write_enable_data_log_force[5443] <= 1'h0;
      write_enable_data_log_force[5444] <= 1'h0;
      write_enable_data_log_force[5445] <= 1'h0;
      write_enable_data_log_force[5446] <= 1'h0;
      write_enable_data_log_force[5447] <= 1'h0;
      write_enable_data_log_force[5448] <= 1'h0;
      write_enable_data_log_force[5449] <= 1'h0;
      write_enable_data_log_force[5450] <= 1'h0;
      write_enable_data_log_force[5451] <= 1'h0;
      write_enable_data_log_force[5452] <= 1'h0;
      write_enable_data_log_force[5453] <= 1'h0;
      write_enable_data_log_force[5454] <= 1'h0;
      write_enable_data_log_force[5455] <= 1'h0;
      write_enable_data_log_force[5456] <= 1'h0;
      write_enable_data_log_force[5457] <= 1'h0;
      write_enable_data_log_force[5458] <= 1'h0;
      write_enable_data_log_force[5459] <= 1'h0;
      write_enable_data_log_force[5460] <= 1'h0;
      write_enable_data_log_force[5461] <= 1'h0;
      write_enable_data_log_force[5462] <= 1'h0;
      write_enable_data_log_force[5463] <= 1'h0;
      write_enable_data_log_force[5464] <= 1'h0;
      write_enable_data_log_force[5465] <= 1'h0;
      write_enable_data_log_force[5466] <= 1'h0;
      write_enable_data_log_force[5467] <= 1'h0;
      write_enable_data_log_force[5468] <= 1'h0;
      write_enable_data_log_force[5469] <= 1'h0;
      write_enable_data_log_force[5470] <= 1'h0;
      write_enable_data_log_force[5471] <= 1'h0;
      write_enable_data_log_force[5472] <= 1'h0;
      write_enable_data_log_force[5473] <= 1'h0;
      write_enable_data_log_force[5474] <= 1'h0;
      write_enable_data_log_force[5475] <= 1'h0;
      write_enable_data_log_force[5476] <= 1'h0;
      write_enable_data_log_force[5477] <= 1'h0;
      write_enable_data_log_force[5478] <= 1'h0;
      write_enable_data_log_force[5479] <= 1'h0;
      write_enable_data_log_force[5480] <= 1'h0;
      write_enable_data_log_force[5481] <= 1'h0;
      write_enable_data_log_force[5482] <= 1'h0;
      write_enable_data_log_force[5483] <= 1'h0;
      write_enable_data_log_force[5484] <= 1'h0;
      write_enable_data_log_force[5485] <= 1'h0;
      write_enable_data_log_force[5486] <= 1'h0;
      write_enable_data_log_force[5487] <= 1'h0;
      write_enable_data_log_force[5488] <= 1'h0;
      write_enable_data_log_force[5489] <= 1'h0;
      write_enable_data_log_force[5490] <= 1'h0;
      write_enable_data_log_force[5491] <= 1'h0;
      write_enable_data_log_force[5492] <= 1'h0;
      write_enable_data_log_force[5493] <= 1'h0;
      write_enable_data_log_force[5494] <= 1'h0;
      write_enable_data_log_force[5495] <= 1'h0;
      write_enable_data_log_force[5496] <= 1'h0;
      write_enable_data_log_force[5497] <= 1'h0;
      write_enable_data_log_force[5498] <= 1'h0;
      write_enable_data_log_force[5499] <= 1'h0;
      write_enable_data_log_force[5500] <= 1'h0;
      write_enable_data_log_force[5501] <= 1'h0;
      write_enable_data_log_force[5502] <= 1'h0;
      write_enable_data_log_force[5503] <= 1'h0;
      write_enable_data_log_force[5504] <= 1'h0;
      write_enable_data_log_force[5505] <= 1'h0;
      write_enable_data_log_force[5506] <= 1'h0;
      write_enable_data_log_force[5507] <= 1'h0;
      write_enable_data_log_force[5508] <= 1'h0;
      write_enable_data_log_force[5509] <= 1'h0;
      write_enable_data_log_force[5510] <= 1'h0;
      write_enable_data_log_force[5511] <= 1'h0;
      write_enable_data_log_force[5512] <= 1'h0;
      write_enable_data_log_force[5513] <= 1'h0;
      write_enable_data_log_force[5514] <= 1'h0;
      write_enable_data_log_force[5515] <= 1'h0;
      write_enable_data_log_force[5516] <= 1'h0;
      write_enable_data_log_force[5517] <= 1'h0;
      write_enable_data_log_force[5518] <= 1'h0;
      write_enable_data_log_force[5519] <= 1'h0;
      write_enable_data_log_force[5520] <= 1'h0;
      write_enable_data_log_force[5521] <= 1'h0;
      write_enable_data_log_force[5522] <= 1'h0;
      write_enable_data_log_force[5523] <= 1'h0;
      write_enable_data_log_force[5524] <= 1'h0;
      write_enable_data_log_force[5525] <= 1'h0;
      write_enable_data_log_force[5526] <= 1'h0;
      write_enable_data_log_force[5527] <= 1'h0;
      write_enable_data_log_force[5528] <= 1'h0;
      write_enable_data_log_force[5529] <= 1'h0;
      write_enable_data_log_force[5530] <= 1'h0;
      write_enable_data_log_force[5531] <= 1'h0;
      write_enable_data_log_force[5532] <= 1'h0;
      write_enable_data_log_force[5533] <= 1'h0;
      write_enable_data_log_force[5534] <= 1'h0;
      write_enable_data_log_force[5535] <= 1'h0;
      write_enable_data_log_force[5536] <= 1'h0;
      write_enable_data_log_force[5537] <= 1'h0;
      write_enable_data_log_force[5538] <= 1'h0;
      write_enable_data_log_force[5539] <= 1'h0;
      write_enable_data_log_force[5540] <= 1'h0;
      write_enable_data_log_force[5541] <= 1'h0;
      write_enable_data_log_force[5542] <= 1'h0;
      write_enable_data_log_force[5543] <= 1'h0;
      write_enable_data_log_force[5544] <= 1'h0;
      write_enable_data_log_force[5545] <= 1'h0;
      write_enable_data_log_force[5546] <= 1'h0;
      write_enable_data_log_force[5547] <= 1'h0;
      write_enable_data_log_force[5548] <= 1'h0;
      write_enable_data_log_force[5549] <= 1'h0;
      write_enable_data_log_force[5550] <= 1'h0;
      write_enable_data_log_force[5551] <= 1'h0;
      write_enable_data_log_force[5552] <= 1'h0;
      write_enable_data_log_force[5553] <= 1'h0;
      write_enable_data_log_force[5554] <= 1'h0;
      write_enable_data_log_force[5555] <= 1'h0;
      write_enable_data_log_force[5556] <= 1'h0;
      write_enable_data_log_force[5557] <= 1'h0;
      write_enable_data_log_force[5558] <= 1'h0;
      write_enable_data_log_force[5559] <= 1'h0;
      write_enable_data_log_force[5560] <= 1'h0;
      write_enable_data_log_force[5561] <= 1'h0;
      write_enable_data_log_force[5562] <= 1'h0;
      write_enable_data_log_force[5563] <= 1'h0;
      write_enable_data_log_force[5564] <= 1'h0;
      write_enable_data_log_force[5565] <= 1'h0;
      write_enable_data_log_force[5566] <= 1'h0;
      write_enable_data_log_force[5567] <= 1'h0;
      write_enable_data_log_force[5568] <= 1'h0;
      write_enable_data_log_force[5569] <= 1'h0;
      write_enable_data_log_force[5570] <= 1'h0;
      write_enable_data_log_force[5571] <= 1'h0;
      write_enable_data_log_force[5572] <= 1'h0;
      write_enable_data_log_force[5573] <= 1'h0;
      write_enable_data_log_force[5574] <= 1'h0;
      write_enable_data_log_force[5575] <= 1'h0;
      write_enable_data_log_force[5576] <= 1'h0;
      write_enable_data_log_force[5577] <= 1'h0;
      write_enable_data_log_force[5578] <= 1'h0;
      write_enable_data_log_force[5579] <= 1'h0;
      write_enable_data_log_force[5580] <= 1'h0;
      write_enable_data_log_force[5581] <= 1'h0;
      write_enable_data_log_force[5582] <= 1'h0;
      write_enable_data_log_force[5583] <= 1'h0;
      write_enable_data_log_force[5584] <= 1'h0;
      write_enable_data_log_force[5585] <= 1'h0;
      write_enable_data_log_force[5586] <= 1'h0;
      write_enable_data_log_force[5587] <= 1'h0;
      write_enable_data_log_force[5588] <= 1'h0;
      write_enable_data_log_force[5589] <= 1'h0;
      write_enable_data_log_force[5590] <= 1'h0;
      write_enable_data_log_force[5591] <= 1'h0;
      write_enable_data_log_force[5592] <= 1'h0;
      write_enable_data_log_force[5593] <= 1'h0;
      write_enable_data_log_force[5594] <= 1'h0;
      write_enable_data_log_force[5595] <= 1'h0;
      write_enable_data_log_force[5596] <= 1'h0;
      write_enable_data_log_force[5597] <= 1'h0;
      write_enable_data_log_force[5598] <= 1'h0;
      write_enable_data_log_force[5599] <= 1'h0;
      write_enable_data_log_force[5600] <= 1'h0;
      write_enable_data_log_force[5601] <= 1'h0;
      write_enable_data_log_force[5602] <= 1'h0;
      write_enable_data_log_force[5603] <= 1'h0;
      write_enable_data_log_force[5604] <= 1'h0;
      write_enable_data_log_force[5605] <= 1'h0;
      write_enable_data_log_force[5606] <= 1'h0;
      write_enable_data_log_force[5607] <= 1'h0;
      write_enable_data_log_force[5608] <= 1'h0;
      write_enable_data_log_force[5609] <= 1'h0;
      write_enable_data_log_force[5610] <= 1'h0;
      write_enable_data_log_force[5611] <= 1'h0;
      write_enable_data_log_force[5612] <= 1'h0;
      write_enable_data_log_force[5613] <= 1'h0;
      write_enable_data_log_force[5614] <= 1'h0;
      write_enable_data_log_force[5615] <= 1'h0;
      write_enable_data_log_force[5616] <= 1'h0;
      write_enable_data_log_force[5617] <= 1'h0;
      write_enable_data_log_force[5618] <= 1'h0;
      write_enable_data_log_force[5619] <= 1'h0;
      write_enable_data_log_force[5620] <= 1'h0;
      write_enable_data_log_force[5621] <= 1'h0;
      write_enable_data_log_force[5622] <= 1'h0;
      write_enable_data_log_force[5623] <= 1'h0;
      write_enable_data_log_force[5624] <= 1'h0;
      write_enable_data_log_force[5625] <= 1'h0;
      write_enable_data_log_force[5626] <= 1'h0;
      write_enable_data_log_force[5627] <= 1'h0;
      write_enable_data_log_force[5628] <= 1'h0;
      write_enable_data_log_force[5629] <= 1'h0;
      write_enable_data_log_force[5630] <= 1'h0;
      write_enable_data_log_force[5631] <= 1'h0;
      write_enable_data_log_force[5632] <= 1'h0;
      write_enable_data_log_force[5633] <= 1'h0;
      write_enable_data_log_force[5634] <= 1'h0;
      write_enable_data_log_force[5635] <= 1'h0;
      write_enable_data_log_force[5636] <= 1'h0;
      write_enable_data_log_force[5637] <= 1'h0;
      write_enable_data_log_force[5638] <= 1'h0;
      write_enable_data_log_force[5639] <= 1'h0;
      write_enable_data_log_force[5640] <= 1'h0;
      write_enable_data_log_force[5641] <= 1'h0;
      write_enable_data_log_force[5642] <= 1'h0;
      write_enable_data_log_force[5643] <= 1'h0;
      write_enable_data_log_force[5644] <= 1'h0;
      write_enable_data_log_force[5645] <= 1'h0;
      write_enable_data_log_force[5646] <= 1'h0;
      write_enable_data_log_force[5647] <= 1'h0;
      write_enable_data_log_force[5648] <= 1'h0;
      write_enable_data_log_force[5649] <= 1'h0;
      write_enable_data_log_force[5650] <= 1'h0;
      write_enable_data_log_force[5651] <= 1'h0;
      write_enable_data_log_force[5652] <= 1'h0;
      write_enable_data_log_force[5653] <= 1'h0;
      write_enable_data_log_force[5654] <= 1'h0;
      write_enable_data_log_force[5655] <= 1'h0;
      write_enable_data_log_force[5656] <= 1'h0;
      write_enable_data_log_force[5657] <= 1'h0;
      write_enable_data_log_force[5658] <= 1'h0;
      write_enable_data_log_force[5659] <= 1'h0;
      write_enable_data_log_force[5660] <= 1'h0;
      write_enable_data_log_force[5661] <= 1'h0;
      write_enable_data_log_force[5662] <= 1'h0;
      write_enable_data_log_force[5663] <= 1'h0;
      write_enable_data_log_force[5664] <= 1'h0;
      write_enable_data_log_force[5665] <= 1'h0;
      write_enable_data_log_force[5666] <= 1'h0;
      write_enable_data_log_force[5667] <= 1'h0;
      write_enable_data_log_force[5668] <= 1'h0;
      write_enable_data_log_force[5669] <= 1'h0;
      write_enable_data_log_force[5670] <= 1'h0;
      write_enable_data_log_force[5671] <= 1'h0;
      write_enable_data_log_force[5672] <= 1'h0;
      write_enable_data_log_force[5673] <= 1'h0;
      write_enable_data_log_force[5674] <= 1'h0;
      write_enable_data_log_force[5675] <= 1'h0;
      write_enable_data_log_force[5676] <= 1'h0;
      write_enable_data_log_force[5677] <= 1'h0;
      write_enable_data_log_force[5678] <= 1'h0;
      write_enable_data_log_force[5679] <= 1'h0;
      write_enable_data_log_force[5680] <= 1'h0;
      write_enable_data_log_force[5681] <= 1'h0;
      write_enable_data_log_force[5682] <= 1'h0;
      write_enable_data_log_force[5683] <= 1'h0;
      write_enable_data_log_force[5684] <= 1'h0;
      write_enable_data_log_force[5685] <= 1'h0;
      write_enable_data_log_force[5686] <= 1'h0;
      write_enable_data_log_force[5687] <= 1'h0;
      write_enable_data_log_force[5688] <= 1'h0;
      write_enable_data_log_force[5689] <= 1'h0;
      write_enable_data_log_force[5690] <= 1'h0;
      write_enable_data_log_force[5691] <= 1'h0;
      write_enable_data_log_force[5692] <= 1'h0;
      write_enable_data_log_force[5693] <= 1'h0;
      write_enable_data_log_force[5694] <= 1'h0;
      write_enable_data_log_force[5695] <= 1'h0;
      write_enable_data_log_force[5696] <= 1'h0;
      write_enable_data_log_force[5697] <= 1'h0;
      write_enable_data_log_force[5698] <= 1'h0;
      write_enable_data_log_force[5699] <= 1'h0;
      write_enable_data_log_force[5700] <= 1'h0;
      write_enable_data_log_force[5701] <= 1'h0;
      write_enable_data_log_force[5702] <= 1'h0;
      write_enable_data_log_force[5703] <= 1'h0;
      write_enable_data_log_force[5704] <= 1'h0;
      write_enable_data_log_force[5705] <= 1'h0;
      write_enable_data_log_force[5706] <= 1'h0;
      write_enable_data_log_force[5707] <= 1'h0;
      write_enable_data_log_force[5708] <= 1'h0;
      write_enable_data_log_force[5709] <= 1'h0;
      write_enable_data_log_force[5710] <= 1'h0;
      write_enable_data_log_force[5711] <= 1'h0;
      write_enable_data_log_force[5712] <= 1'h0;
      write_enable_data_log_force[5713] <= 1'h0;
      write_enable_data_log_force[5714] <= 1'h0;
      write_enable_data_log_force[5715] <= 1'h0;
      write_enable_data_log_force[5716] <= 1'h0;
      write_enable_data_log_force[5717] <= 1'h0;
      write_enable_data_log_force[5718] <= 1'h0;
      write_enable_data_log_force[5719] <= 1'h0;
      write_enable_data_log_force[5720] <= 1'h0;
      write_enable_data_log_force[5721] <= 1'h0;
      write_enable_data_log_force[5722] <= 1'h0;
      write_enable_data_log_force[5723] <= 1'h0;
      write_enable_data_log_force[5724] <= 1'h0;
      write_enable_data_log_force[5725] <= 1'h0;
      write_enable_data_log_force[5726] <= 1'h0;
      write_enable_data_log_force[5727] <= 1'h0;
      write_enable_data_log_force[5728] <= 1'h0;
      write_enable_data_log_force[5729] <= 1'h0;
      write_enable_data_log_force[5730] <= 1'h0;
      write_enable_data_log_force[5731] <= 1'h0;
      write_enable_data_log_force[5732] <= 1'h0;
      write_enable_data_log_force[5733] <= 1'h0;
      write_enable_data_log_force[5734] <= 1'h0;
      write_enable_data_log_force[5735] <= 1'h0;
      write_enable_data_log_force[5736] <= 1'h0;
      write_enable_data_log_force[5737] <= 1'h0;
      write_enable_data_log_force[5738] <= 1'h0;
      write_enable_data_log_force[5739] <= 1'h0;
      write_enable_data_log_force[5740] <= 1'h0;
      write_enable_data_log_force[5741] <= 1'h0;
      write_enable_data_log_force[5742] <= 1'h0;
      write_enable_data_log_force[5743] <= 1'h0;
      write_enable_data_log_force[5744] <= 1'h0;
      write_enable_data_log_force[5745] <= 1'h0;
      write_enable_data_log_force[5746] <= 1'h0;
      write_enable_data_log_force[5747] <= 1'h0;
      write_enable_data_log_force[5748] <= 1'h0;
      write_enable_data_log_force[5749] <= 1'h0;
      write_enable_data_log_force[5750] <= 1'h0;
      write_enable_data_log_force[5751] <= 1'h0;
      write_enable_data_log_force[5752] <= 1'h0;
      write_enable_data_log_force[5753] <= 1'h0;
      write_enable_data_log_force[5754] <= 1'h0;
      write_enable_data_log_force[5755] <= 1'h0;
      write_enable_data_log_force[5756] <= 1'h0;
      write_enable_data_log_force[5757] <= 1'h0;
      write_enable_data_log_force[5758] <= 1'h0;
      write_enable_data_log_force[5759] <= 1'h0;
      write_enable_data_log_force[5760] <= 1'h0;
      write_enable_data_log_force[5761] <= 1'h0;
      write_enable_data_log_force[5762] <= 1'h0;
      write_enable_data_log_force[5763] <= 1'h0;
      write_enable_data_log_force[5764] <= 1'h0;
      write_enable_data_log_force[5765] <= 1'h0;
      write_enable_data_log_force[5766] <= 1'h0;
      write_enable_data_log_force[5767] <= 1'h0;
      write_enable_data_log_force[5768] <= 1'h0;
      write_enable_data_log_force[5769] <= 1'h0;
      write_enable_data_log_force[5770] <= 1'h0;
      write_enable_data_log_force[5771] <= 1'h0;
      write_enable_data_log_force[5772] <= 1'h0;
      write_enable_data_log_force[5773] <= 1'h0;
      write_enable_data_log_force[5774] <= 1'h0;
      write_enable_data_log_force[5775] <= 1'h0;
      write_enable_data_log_force[5776] <= 1'h0;
      write_enable_data_log_force[5777] <= 1'h0;
      write_enable_data_log_force[5778] <= 1'h0;
      write_enable_data_log_force[5779] <= 1'h0;
      write_enable_data_log_force[5780] <= 1'h0;
      write_enable_data_log_force[5781] <= 1'h0;
      write_enable_data_log_force[5782] <= 1'h0;
      write_enable_data_log_force[5783] <= 1'h0;
      write_enable_data_log_force[5784] <= 1'h0;
      write_enable_data_log_force[5785] <= 1'h0;
      write_enable_data_log_force[5786] <= 1'h0;
      write_enable_data_log_force[5787] <= 1'h0;
      write_enable_data_log_force[5788] <= 1'h0;
      write_enable_data_log_force[5789] <= 1'h0;
      write_enable_data_log_force[5790] <= 1'h0;
      write_enable_data_log_force[5791] <= 1'h0;
      write_enable_data_log_force[5792] <= 1'h0;
      write_enable_data_log_force[5793] <= 1'h0;
      write_enable_data_log_force[5794] <= 1'h0;
      write_enable_data_log_force[5795] <= 1'h0;
      write_enable_data_log_force[5796] <= 1'h0;
      write_enable_data_log_force[5797] <= 1'h0;
      write_enable_data_log_force[5798] <= 1'h0;
      write_enable_data_log_force[5799] <= 1'h0;
      write_enable_data_log_force[5800] <= 1'h0;
      write_enable_data_log_force[5801] <= 1'h0;
      write_enable_data_log_force[5802] <= 1'h0;
      write_enable_data_log_force[5803] <= 1'h0;
      write_enable_data_log_force[5804] <= 1'h0;
      write_enable_data_log_force[5805] <= 1'h0;
      write_enable_data_log_force[5806] <= 1'h0;
      write_enable_data_log_force[5807] <= 1'h0;
      write_enable_data_log_force[5808] <= 1'h0;
      write_enable_data_log_force[5809] <= 1'h0;
      write_enable_data_log_force[5810] <= 1'h0;
      write_enable_data_log_force[5811] <= 1'h0;
      write_enable_data_log_force[5812] <= 1'h0;
      write_enable_data_log_force[5813] <= 1'h0;
      write_enable_data_log_force[5814] <= 1'h0;
      write_enable_data_log_force[5815] <= 1'h0;
      write_enable_data_log_force[5816] <= 1'h0;
      write_enable_data_log_force[5817] <= 1'h0;
      write_enable_data_log_force[5818] <= 1'h0;
      write_enable_data_log_force[5819] <= 1'h0;
      write_enable_data_log_force[5820] <= 1'h0;
      write_enable_data_log_force[5821] <= 1'h0;
      write_enable_data_log_force[5822] <= 1'h0;
      write_enable_data_log_force[5823] <= 1'h0;
      write_enable_data_log_force[5824] <= 1'h0;
      write_enable_data_log_force[5825] <= 1'h0;
      write_enable_data_log_force[5826] <= 1'h0;
      write_enable_data_log_force[5827] <= 1'h0;
      write_enable_data_log_force[5828] <= 1'h0;
      write_enable_data_log_force[5829] <= 1'h0;
      write_enable_data_log_force[5830] <= 1'h0;
      write_enable_data_log_force[5831] <= 1'h0;
      write_enable_data_log_force[5832] <= 1'h0;
      write_enable_data_log_force[5833] <= 1'h0;
      write_enable_data_log_force[5834] <= 1'h0;
      write_enable_data_log_force[5835] <= 1'h0;
      write_enable_data_log_force[5836] <= 1'h0;
      write_enable_data_log_force[5837] <= 1'h0;
      write_enable_data_log_force[5838] <= 1'h0;
      write_enable_data_log_force[5839] <= 1'h0;
      write_enable_data_log_force[5840] <= 1'h0;
      write_enable_data_log_force[5841] <= 1'h0;
      write_enable_data_log_force[5842] <= 1'h0;
      write_enable_data_log_force[5843] <= 1'h0;
      write_enable_data_log_force[5844] <= 1'h0;
      write_enable_data_log_force[5845] <= 1'h0;
      write_enable_data_log_force[5846] <= 1'h0;
      write_enable_data_log_force[5847] <= 1'h0;
      write_enable_data_log_force[5848] <= 1'h0;
      write_enable_data_log_force[5849] <= 1'h0;
      write_enable_data_log_force[5850] <= 1'h0;
      write_enable_data_log_force[5851] <= 1'h0;
      write_enable_data_log_force[5852] <= 1'h0;
      write_enable_data_log_force[5853] <= 1'h0;
      write_enable_data_log_force[5854] <= 1'h0;
      write_enable_data_log_force[5855] <= 1'h0;
      write_enable_data_log_force[5856] <= 1'h0;
      write_enable_data_log_force[5857] <= 1'h0;
      write_enable_data_log_force[5858] <= 1'h0;
      write_enable_data_log_force[5859] <= 1'h0;
      write_enable_data_log_force[5860] <= 1'h0;
      write_enable_data_log_force[5861] <= 1'h0;
      write_enable_data_log_force[5862] <= 1'h0;
      write_enable_data_log_force[5863] <= 1'h0;
      write_enable_data_log_force[5864] <= 1'h0;
      write_enable_data_log_force[5865] <= 1'h0;
      write_enable_data_log_force[5866] <= 1'h0;
      write_enable_data_log_force[5867] <= 1'h0;
      write_enable_data_log_force[5868] <= 1'h0;
      write_enable_data_log_force[5869] <= 1'h0;
      write_enable_data_log_force[5870] <= 1'h0;
      write_enable_data_log_force[5871] <= 1'h0;
      write_enable_data_log_force[5872] <= 1'h0;
      write_enable_data_log_force[5873] <= 1'h0;
      write_enable_data_log_force[5874] <= 1'h0;
      write_enable_data_log_force[5875] <= 1'h0;
      write_enable_data_log_force[5876] <= 1'h0;
      write_enable_data_log_force[5877] <= 1'h0;
      write_enable_data_log_force[5878] <= 1'h0;
      write_enable_data_log_force[5879] <= 1'h0;
      write_enable_data_log_force[5880] <= 1'h0;
      write_enable_data_log_force[5881] <= 1'h0;
      write_enable_data_log_force[5882] <= 1'h0;
      write_enable_data_log_force[5883] <= 1'h0;
      write_enable_data_log_force[5884] <= 1'h0;
      write_enable_data_log_force[5885] <= 1'h0;
      write_enable_data_log_force[5886] <= 1'h0;
      write_enable_data_log_force[5887] <= 1'h0;
      write_enable_data_log_force[5888] <= 1'h0;
      write_enable_data_log_force[5889] <= 1'h0;
      write_enable_data_log_force[5890] <= 1'h0;
      write_enable_data_log_force[5891] <= 1'h0;
      write_enable_data_log_force[5892] <= 1'h0;
      write_enable_data_log_force[5893] <= 1'h0;
      write_enable_data_log_force[5894] <= 1'h0;
      write_enable_data_log_force[5895] <= 1'h0;
      write_enable_data_log_force[5896] <= 1'h0;
      write_enable_data_log_force[5897] <= 1'h0;
      write_enable_data_log_force[5898] <= 1'h0;
      write_enable_data_log_force[5899] <= 1'h0;
      write_enable_data_log_force[5900] <= 1'h0;
      write_enable_data_log_force[5901] <= 1'h0;
      write_enable_data_log_force[5902] <= 1'h0;
      write_enable_data_log_force[5903] <= 1'h0;
      write_enable_data_log_force[5904] <= 1'h0;
      write_enable_data_log_force[5905] <= 1'h0;
      write_enable_data_log_force[5906] <= 1'h0;
      write_enable_data_log_force[5907] <= 1'h0;
      write_enable_data_log_force[5908] <= 1'h0;
      write_enable_data_log_force[5909] <= 1'h0;
      write_enable_data_log_force[5910] <= 1'h0;
      write_enable_data_log_force[5911] <= 1'h0;
      write_enable_data_log_force[5912] <= 1'h0;
      write_enable_data_log_force[5913] <= 1'h0;
      write_enable_data_log_force[5914] <= 1'h0;
      write_enable_data_log_force[5915] <= 1'h0;
      write_enable_data_log_force[5916] <= 1'h0;
      write_enable_data_log_force[5917] <= 1'h0;
      write_enable_data_log_force[5918] <= 1'h0;
      write_enable_data_log_force[5919] <= 1'h0;
      write_enable_data_log_force[5920] <= 1'h0;
      write_enable_data_log_force[5921] <= 1'h0;
      write_enable_data_log_force[5922] <= 1'h0;
      write_enable_data_log_force[5923] <= 1'h0;
      write_enable_data_log_force[5924] <= 1'h0;
      write_enable_data_log_force[5925] <= 1'h0;
      write_enable_data_log_force[5926] <= 1'h0;
      write_enable_data_log_force[5927] <= 1'h0;
      write_enable_data_log_force[5928] <= 1'h0;
      write_enable_data_log_force[5929] <= 1'h0;
      write_enable_data_log_force[5930] <= 1'h0;
      write_enable_data_log_force[5931] <= 1'h0;
      write_enable_data_log_force[5932] <= 1'h0;
      write_enable_data_log_force[5933] <= 1'h0;
      write_enable_data_log_force[5934] <= 1'h0;
      write_enable_data_log_force[5935] <= 1'h0;
      write_enable_data_log_force[5936] <= 1'h0;
      write_enable_data_log_force[5937] <= 1'h0;
      write_enable_data_log_force[5938] <= 1'h0;
      write_enable_data_log_force[5939] <= 1'h0;
      write_enable_data_log_force[5940] <= 1'h0;
      write_enable_data_log_force[5941] <= 1'h0;
      write_enable_data_log_force[5942] <= 1'h0;
      write_enable_data_log_force[5943] <= 1'h0;
      write_enable_data_log_force[5944] <= 1'h0;
      write_enable_data_log_force[5945] <= 1'h0;
      write_enable_data_log_force[5946] <= 1'h0;
      write_enable_data_log_force[5947] <= 1'h0;
      write_enable_data_log_force[5948] <= 1'h0;
      write_enable_data_log_force[5949] <= 1'h0;
      write_enable_data_log_force[5950] <= 1'h0;
      write_enable_data_log_force[5951] <= 1'h0;
      write_enable_data_log_force[5952] <= 1'h0;
      write_enable_data_log_force[5953] <= 1'h0;
      write_enable_data_log_force[5954] <= 1'h0;
      write_enable_data_log_force[5955] <= 1'h0;
      write_enable_data_log_force[5956] <= 1'h0;
      write_enable_data_log_force[5957] <= 1'h0;
      write_enable_data_log_force[5958] <= 1'h0;
      write_enable_data_log_force[5959] <= 1'h0;
      write_enable_data_log_force[5960] <= 1'h0;
      write_enable_data_log_force[5961] <= 1'h0;
      write_enable_data_log_force[5962] <= 1'h0;
      write_enable_data_log_force[5963] <= 1'h0;
      write_enable_data_log_force[5964] <= 1'h0;
      write_enable_data_log_force[5965] <= 1'h0;
      write_enable_data_log_force[5966] <= 1'h0;
      write_enable_data_log_force[5967] <= 1'h0;
      write_enable_data_log_force[5968] <= 1'h0;
      write_enable_data_log_force[5969] <= 1'h0;
      write_enable_data_log_force[5970] <= 1'h0;
      write_enable_data_log_force[5971] <= 1'h0;
      write_enable_data_log_force[5972] <= 1'h0;
      write_enable_data_log_force[5973] <= 1'h0;
      write_enable_data_log_force[5974] <= 1'h0;
      write_enable_data_log_force[5975] <= 1'h0;
      write_enable_data_log_force[5976] <= 1'h0;
      write_enable_data_log_force[5977] <= 1'h0;
      write_enable_data_log_force[5978] <= 1'h0;
      write_enable_data_log_force[5979] <= 1'h0;
      write_enable_data_log_force[5980] <= 1'h0;
      write_enable_data_log_force[5981] <= 1'h0;
      write_enable_data_log_force[5982] <= 1'h0;
      write_enable_data_log_force[5983] <= 1'h0;
      write_enable_data_log_force[5984] <= 1'h0;
      write_enable_data_log_force[5985] <= 1'h0;
      write_enable_data_log_force[5986] <= 1'h0;
      write_enable_data_log_force[5987] <= 1'h0;
      write_enable_data_log_force[5988] <= 1'h0;
      write_enable_data_log_force[5989] <= 1'h0;
      write_enable_data_log_force[5990] <= 1'h0;
      write_enable_data_log_force[5991] <= 1'h0;
      write_enable_data_log_force[5992] <= 1'h0;
      write_enable_data_log_force[5993] <= 1'h0;
      write_enable_data_log_force[5994] <= 1'h0;
      write_enable_data_log_force[5995] <= 1'h0;
      write_enable_data_log_force[5996] <= 1'h0;
      write_enable_data_log_force[5997] <= 1'h0;
      write_enable_data_log_force[5998] <= 1'h0;
      write_enable_data_log_force[5999] <= 1'h0;
      write_enable_data_log_force[6000] <= 1'h0;
      write_enable_data_log_force[6001] <= 1'h0;
      write_enable_data_log_force[6002] <= 1'h0;
      write_enable_data_log_force[6003] <= 1'h0;
      write_enable_data_log_force[6004] <= 1'h0;
      write_enable_data_log_force[6005] <= 1'h0;
      write_enable_data_log_force[6006] <= 1'h0;
      write_enable_data_log_force[6007] <= 1'h0;
      write_enable_data_log_force[6008] <= 1'h0;
      write_enable_data_log_force[6009] <= 1'h0;
      write_enable_data_log_force[6010] <= 1'h0;
      write_enable_data_log_force[6011] <= 1'h0;
      write_enable_data_log_force[6012] <= 1'h0;
      write_enable_data_log_force[6013] <= 1'h0;
      write_enable_data_log_force[6014] <= 1'h0;
      write_enable_data_log_force[6015] <= 1'h0;
      write_enable_data_log_force[6016] <= 1'h0;
      write_enable_data_log_force[6017] <= 1'h0;
      write_enable_data_log_force[6018] <= 1'h0;
      write_enable_data_log_force[6019] <= 1'h0;
      write_enable_data_log_force[6020] <= 1'h0;
      write_enable_data_log_force[6021] <= 1'h0;
      write_enable_data_log_force[6022] <= 1'h0;
      write_enable_data_log_force[6023] <= 1'h0;
      write_enable_data_log_force[6024] <= 1'h0;
      write_enable_data_log_force[6025] <= 1'h0;
      write_enable_data_log_force[6026] <= 1'h0;
      write_enable_data_log_force[6027] <= 1'h0;
      write_enable_data_log_force[6028] <= 1'h0;
      write_enable_data_log_force[6029] <= 1'h0;
      write_enable_data_log_force[6030] <= 1'h0;
      write_enable_data_log_force[6031] <= 1'h0;
      write_enable_data_log_force[6032] <= 1'h0;
      write_enable_data_log_force[6033] <= 1'h0;
      write_enable_data_log_force[6034] <= 1'h0;
      write_enable_data_log_force[6035] <= 1'h0;
      write_enable_data_log_force[6036] <= 1'h0;
      write_enable_data_log_force[6037] <= 1'h0;
      write_enable_data_log_force[6038] <= 1'h0;
      write_enable_data_log_force[6039] <= 1'h0;
      write_enable_data_log_force[6040] <= 1'h0;
      write_enable_data_log_force[6041] <= 1'h0;
      write_enable_data_log_force[6042] <= 1'h0;
      write_enable_data_log_force[6043] <= 1'h0;
      write_enable_data_log_force[6044] <= 1'h0;
      write_enable_data_log_force[6045] <= 1'h0;
      write_enable_data_log_force[6046] <= 1'h0;
      write_enable_data_log_force[6047] <= 1'h0;
      write_enable_data_log_force[6048] <= 1'h0;
      write_enable_data_log_force[6049] <= 1'h0;
      write_enable_data_log_force[6050] <= 1'h0;
      write_enable_data_log_force[6051] <= 1'h0;
      write_enable_data_log_force[6052] <= 1'h0;
      write_enable_data_log_force[6053] <= 1'h0;
      write_enable_data_log_force[6054] <= 1'h0;
      write_enable_data_log_force[6055] <= 1'h0;
      write_enable_data_log_force[6056] <= 1'h0;
      write_enable_data_log_force[6057] <= 1'h0;
      write_enable_data_log_force[6058] <= 1'h0;
      write_enable_data_log_force[6059] <= 1'h0;
      write_enable_data_log_force[6060] <= 1'h0;
      write_enable_data_log_force[6061] <= 1'h0;
      write_enable_data_log_force[6062] <= 1'h0;
      write_enable_data_log_force[6063] <= 1'h0;
      write_enable_data_log_force[6064] <= 1'h0;
      write_enable_data_log_force[6065] <= 1'h0;
      write_enable_data_log_force[6066] <= 1'h0;
      write_enable_data_log_force[6067] <= 1'h0;
      write_enable_data_log_force[6068] <= 1'h0;
      write_enable_data_log_force[6069] <= 1'h0;
      write_enable_data_log_force[6070] <= 1'h0;
      write_enable_data_log_force[6071] <= 1'h0;
      write_enable_data_log_force[6072] <= 1'h0;
      write_enable_data_log_force[6073] <= 1'h0;
      write_enable_data_log_force[6074] <= 1'h0;
      write_enable_data_log_force[6075] <= 1'h0;
      write_enable_data_log_force[6076] <= 1'h0;
      write_enable_data_log_force[6077] <= 1'h0;
      write_enable_data_log_force[6078] <= 1'h0;
      write_enable_data_log_force[6079] <= 1'h0;
      write_enable_data_log_force[6080] <= 1'h0;
      write_enable_data_log_force[6081] <= 1'h0;
      write_enable_data_log_force[6082] <= 1'h0;
      write_enable_data_log_force[6083] <= 1'h0;
      write_enable_data_log_force[6084] <= 1'h0;
      write_enable_data_log_force[6085] <= 1'h0;
      write_enable_data_log_force[6086] <= 1'h0;
      write_enable_data_log_force[6087] <= 1'h0;
      write_enable_data_log_force[6088] <= 1'h0;
      write_enable_data_log_force[6089] <= 1'h0;
      write_enable_data_log_force[6090] <= 1'h0;
      write_enable_data_log_force[6091] <= 1'h0;
      write_enable_data_log_force[6092] <= 1'h0;
      write_enable_data_log_force[6093] <= 1'h0;
      write_enable_data_log_force[6094] <= 1'h0;
      write_enable_data_log_force[6095] <= 1'h0;
      write_enable_data_log_force[6096] <= 1'h0;
      write_enable_data_log_force[6097] <= 1'h0;
      write_enable_data_log_force[6098] <= 1'h0;
      write_enable_data_log_force[6099] <= 1'h0;
      write_enable_data_log_force[6100] <= 1'h0;
      write_enable_data_log_force[6101] <= 1'h0;
      write_enable_data_log_force[6102] <= 1'h0;
      write_enable_data_log_force[6103] <= 1'h0;
      write_enable_data_log_force[6104] <= 1'h0;
      write_enable_data_log_force[6105] <= 1'h0;
      write_enable_data_log_force[6106] <= 1'h0;
      write_enable_data_log_force[6107] <= 1'h0;
      write_enable_data_log_force[6108] <= 1'h0;
      write_enable_data_log_force[6109] <= 1'h0;
      write_enable_data_log_force[6110] <= 1'h0;
      write_enable_data_log_force[6111] <= 1'h0;
      write_enable_data_log_force[6112] <= 1'h0;
      write_enable_data_log_force[6113] <= 1'h0;
      write_enable_data_log_force[6114] <= 1'h0;
      write_enable_data_log_force[6115] <= 1'h0;
      write_enable_data_log_force[6116] <= 1'h0;
      write_enable_data_log_force[6117] <= 1'h0;
      write_enable_data_log_force[6118] <= 1'h0;
      write_enable_data_log_force[6119] <= 1'h0;
      write_enable_data_log_force[6120] <= 1'h0;
      write_enable_data_log_force[6121] <= 1'h0;
      write_enable_data_log_force[6122] <= 1'h0;
      write_enable_data_log_force[6123] <= 1'h0;
      write_enable_data_log_force[6124] <= 1'h0;
      write_enable_data_log_force[6125] <= 1'h0;
      write_enable_data_log_force[6126] <= 1'h0;
      write_enable_data_log_force[6127] <= 1'h0;
      write_enable_data_log_force[6128] <= 1'h0;
      write_enable_data_log_force[6129] <= 1'h0;
      write_enable_data_log_force[6130] <= 1'h0;
      write_enable_data_log_force[6131] <= 1'h0;
      write_enable_data_log_force[6132] <= 1'h0;
      write_enable_data_log_force[6133] <= 1'h0;
      write_enable_data_log_force[6134] <= 1'h0;
      write_enable_data_log_force[6135] <= 1'h0;
      write_enable_data_log_force[6136] <= 1'h0;
      write_enable_data_log_force[6137] <= 1'h0;
      write_enable_data_log_force[6138] <= 1'h0;
      write_enable_data_log_force[6139] <= 1'h0;
      write_enable_data_log_force[6140] <= 1'h0;
      write_enable_data_log_force[6141] <= 1'h0;
      write_enable_data_log_force[6142] <= 1'h0;
      write_enable_data_log_force[6143] <= 1'h0;
      write_enable_data_log_force[6144] <= 1'h0;
      write_enable_data_log_force[6145] <= 1'h0;
      write_enable_data_log_force[6146] <= 1'h0;
      write_enable_data_log_force[6147] <= 1'h0;
      write_enable_data_log_force[6148] <= 1'h0;
      write_enable_data_log_force[6149] <= 1'h0;
      write_enable_data_log_force[6150] <= 1'h0;
      write_enable_data_log_force[6151] <= 1'h0;
      write_enable_data_log_force[6152] <= 1'h0;
      write_enable_data_log_force[6153] <= 1'h0;
      write_enable_data_log_force[6154] <= 1'h0;
      write_enable_data_log_force[6155] <= 1'h0;
      write_enable_data_log_force[6156] <= 1'h0;
      write_enable_data_log_force[6157] <= 1'h0;
      write_enable_data_log_force[6158] <= 1'h0;
      write_enable_data_log_force[6159] <= 1'h0;
      write_enable_data_log_force[6160] <= 1'h0;
      write_enable_data_log_force[6161] <= 1'h0;
      write_enable_data_log_force[6162] <= 1'h0;
      write_enable_data_log_force[6163] <= 1'h0;
      write_enable_data_log_force[6164] <= 1'h0;
      write_enable_data_log_force[6165] <= 1'h0;
      write_enable_data_log_force[6166] <= 1'h0;
      write_enable_data_log_force[6167] <= 1'h0;
      write_enable_data_log_force[6168] <= 1'h0;
      write_enable_data_log_force[6169] <= 1'h0;
      write_enable_data_log_force[6170] <= 1'h0;
      write_enable_data_log_force[6171] <= 1'h0;
      write_enable_data_log_force[6172] <= 1'h0;
      write_enable_data_log_force[6173] <= 1'h0;
      write_enable_data_log_force[6174] <= 1'h0;
      write_enable_data_log_force[6175] <= 1'h0;
      write_enable_data_log_force[6176] <= 1'h0;
      write_enable_data_log_force[6177] <= 1'h0;
      write_enable_data_log_force[6178] <= 1'h0;
      write_enable_data_log_force[6179] <= 1'h0;
      write_enable_data_log_force[6180] <= 1'h0;
      write_enable_data_log_force[6181] <= 1'h0;
      write_enable_data_log_force[6182] <= 1'h0;
      write_enable_data_log_force[6183] <= 1'h0;
      write_enable_data_log_force[6184] <= 1'h0;
      write_enable_data_log_force[6185] <= 1'h0;
      write_enable_data_log_force[6186] <= 1'h0;
      write_enable_data_log_force[6187] <= 1'h0;
      write_enable_data_log_force[6188] <= 1'h0;
      write_enable_data_log_force[6189] <= 1'h0;
      write_enable_data_log_force[6190] <= 1'h0;
      write_enable_data_log_force[6191] <= 1'h0;
      write_enable_data_log_force[6192] <= 1'h0;
      write_enable_data_log_force[6193] <= 1'h0;
      write_enable_data_log_force[6194] <= 1'h0;
      write_enable_data_log_force[6195] <= 1'h0;
      write_enable_data_log_force[6196] <= 1'h0;
      write_enable_data_log_force[6197] <= 1'h0;
      write_enable_data_log_force[6198] <= 1'h0;
      write_enable_data_log_force[6199] <= 1'h0;
      write_enable_data_log_force[6200] <= 1'h0;
      write_enable_data_log_force[6201] <= 1'h0;
      write_enable_data_log_force[6202] <= 1'h0;
      write_enable_data_log_force[6203] <= 1'h0;
      write_enable_data_log_force[6204] <= 1'h0;
      write_enable_data_log_force[6205] <= 1'h0;
      write_enable_data_log_force[6206] <= 1'h0;
      write_enable_data_log_force[6207] <= 1'h0;
      write_enable_data_log_force[6208] <= 1'h0;
      write_enable_data_log_force[6209] <= 1'h0;
      write_enable_data_log_force[6210] <= 1'h0;
      write_enable_data_log_force[6211] <= 1'h0;
      write_enable_data_log_force[6212] <= 1'h0;
      write_enable_data_log_force[6213] <= 1'h0;
      write_enable_data_log_force[6214] <= 1'h0;
      write_enable_data_log_force[6215] <= 1'h0;
      write_enable_data_log_force[6216] <= 1'h0;
      write_enable_data_log_force[6217] <= 1'h0;
      write_enable_data_log_force[6218] <= 1'h0;
      write_enable_data_log_force[6219] <= 1'h0;
      write_enable_data_log_force[6220] <= 1'h0;
      write_enable_data_log_force[6221] <= 1'h0;
      write_enable_data_log_force[6222] <= 1'h0;
      write_enable_data_log_force[6223] <= 1'h0;
      write_enable_data_log_force[6224] <= 1'h0;
      write_enable_data_log_force[6225] <= 1'h0;
      write_enable_data_log_force[6226] <= 1'h0;
      write_enable_data_log_force[6227] <= 1'h0;
      write_enable_data_log_force[6228] <= 1'h0;
      write_enable_data_log_force[6229] <= 1'h0;
      write_enable_data_log_force[6230] <= 1'h0;
      write_enable_data_log_force[6231] <= 1'h0;
      write_enable_data_log_force[6232] <= 1'h0;
      write_enable_data_log_force[6233] <= 1'h0;
      write_enable_data_log_force[6234] <= 1'h0;
      write_enable_data_log_force[6235] <= 1'h0;
      write_enable_data_log_force[6236] <= 1'h0;
      write_enable_data_log_force[6237] <= 1'h0;
      write_enable_data_log_force[6238] <= 1'h0;
      write_enable_data_log_force[6239] <= 1'h0;
      write_enable_data_log_force[6240] <= 1'h0;
      write_enable_data_log_force[6241] <= 1'h0;
      write_enable_data_log_force[6242] <= 1'h0;
      write_enable_data_log_force[6243] <= 1'h0;
      write_enable_data_log_force[6244] <= 1'h0;
      write_enable_data_log_force[6245] <= 1'h0;
      write_enable_data_log_force[6246] <= 1'h0;
      write_enable_data_log_force[6247] <= 1'h0;
      write_enable_data_log_force[6248] <= 1'h0;
      write_enable_data_log_force[6249] <= 1'h0;
      write_enable_data_log_force[6250] <= 1'h0;
      write_enable_data_log_force[6251] <= 1'h0;
      write_enable_data_log_force[6252] <= 1'h0;
      write_enable_data_log_force[6253] <= 1'h0;
      write_enable_data_log_force[6254] <= 1'h0;
      write_enable_data_log_force[6255] <= 1'h0;
      write_enable_data_log_force[6256] <= 1'h0;
      write_enable_data_log_force[6257] <= 1'h0;
      write_enable_data_log_force[6258] <= 1'h0;
      write_enable_data_log_force[6259] <= 1'h0;
      write_enable_data_log_force[6260] <= 1'h0;
      write_enable_data_log_force[6261] <= 1'h0;
      write_enable_data_log_force[6262] <= 1'h0;
      write_enable_data_log_force[6263] <= 1'h0;
      write_enable_data_log_force[6264] <= 1'h0;
      write_enable_data_log_force[6265] <= 1'h0;
      write_enable_data_log_force[6266] <= 1'h0;
      write_enable_data_log_force[6267] <= 1'h0;
      write_enable_data_log_force[6268] <= 1'h0;
      write_enable_data_log_force[6269] <= 1'h0;
      write_enable_data_log_force[6270] <= 1'h0;
      write_enable_data_log_force[6271] <= 1'h0;
      write_enable_data_log_force[6272] <= 1'h0;
      write_enable_data_log_force[6273] <= 1'h0;
      write_enable_data_log_force[6274] <= 1'h0;
      write_enable_data_log_force[6275] <= 1'h0;
      write_enable_data_log_force[6276] <= 1'h0;
      write_enable_data_log_force[6277] <= 1'h0;
      write_enable_data_log_force[6278] <= 1'h0;
      write_enable_data_log_force[6279] <= 1'h0;
      write_enable_data_log_force[6280] <= 1'h0;
      write_enable_data_log_force[6281] <= 1'h0;
      write_enable_data_log_force[6282] <= 1'h0;
      write_enable_data_log_force[6283] <= 1'h0;
      write_enable_data_log_force[6284] <= 1'h0;
      write_enable_data_log_force[6285] <= 1'h0;
      write_enable_data_log_force[6286] <= 1'h0;
      write_enable_data_log_force[6287] <= 1'h0;
      write_enable_data_log_force[6288] <= 1'h0;
      write_enable_data_log_force[6289] <= 1'h0;
      write_enable_data_log_force[6290] <= 1'h0;
      write_enable_data_log_force[6291] <= 1'h0;
      write_enable_data_log_force[6292] <= 1'h0;
      write_enable_data_log_force[6293] <= 1'h0;
      write_enable_data_log_force[6294] <= 1'h0;
      write_enable_data_log_force[6295] <= 1'h0;
      write_enable_data_log_force[6296] <= 1'h0;
      write_enable_data_log_force[6297] <= 1'h0;
      write_enable_data_log_force[6298] <= 1'h0;
      write_enable_data_log_force[6299] <= 1'h0;
      write_enable_data_log_force[6300] <= 1'h0;
      write_enable_data_log_force[6301] <= 1'h0;
      write_enable_data_log_force[6302] <= 1'h0;
      write_enable_data_log_force[6303] <= 1'h0;
      write_enable_data_log_force[6304] <= 1'h0;
      write_enable_data_log_force[6305] <= 1'h0;
      write_enable_data_log_force[6306] <= 1'h0;
      write_enable_data_log_force[6307] <= 1'h0;
      write_enable_data_log_force[6308] <= 1'h0;
      write_enable_data_log_force[6309] <= 1'h0;
      write_enable_data_log_force[6310] <= 1'h0;
      write_enable_data_log_force[6311] <= 1'h0;
      write_enable_data_log_force[6312] <= 1'h0;
      write_enable_data_log_force[6313] <= 1'h0;
      write_enable_data_log_force[6314] <= 1'h0;
      write_enable_data_log_force[6315] <= 1'h0;
      write_enable_data_log_force[6316] <= 1'h0;
      write_enable_data_log_force[6317] <= 1'h0;
      write_enable_data_log_force[6318] <= 1'h0;
      write_enable_data_log_force[6319] <= 1'h0;
      write_enable_data_log_force[6320] <= 1'h0;
      write_enable_data_log_force[6321] <= 1'h0;
      write_enable_data_log_force[6322] <= 1'h0;
      write_enable_data_log_force[6323] <= 1'h0;
      write_enable_data_log_force[6324] <= 1'h0;
      write_enable_data_log_force[6325] <= 1'h0;
      write_enable_data_log_force[6326] <= 1'h0;
      write_enable_data_log_force[6327] <= 1'h0;
      write_enable_data_log_force[6328] <= 1'h0;
      write_enable_data_log_force[6329] <= 1'h0;
      write_enable_data_log_force[6330] <= 1'h0;
      write_enable_data_log_force[6331] <= 1'h0;
      write_enable_data_log_force[6332] <= 1'h0;
      write_enable_data_log_force[6333] <= 1'h0;
      write_enable_data_log_force[6334] <= 1'h0;
      write_enable_data_log_force[6335] <= 1'h0;
      write_enable_data_log_force[6336] <= 1'h0;
      write_enable_data_log_force[6337] <= 1'h0;
      write_enable_data_log_force[6338] <= 1'h0;
      write_enable_data_log_force[6339] <= 1'h0;
      write_enable_data_log_force[6340] <= 1'h0;
      write_enable_data_log_force[6341] <= 1'h0;
      write_enable_data_log_force[6342] <= 1'h0;
      write_enable_data_log_force[6343] <= 1'h0;
      write_enable_data_log_force[6344] <= 1'h0;
      write_enable_data_log_force[6345] <= 1'h0;
      write_enable_data_log_force[6346] <= 1'h0;
      write_enable_data_log_force[6347] <= 1'h0;
      write_enable_data_log_force[6348] <= 1'h0;
      write_enable_data_log_force[6349] <= 1'h0;
      write_enable_data_log_force[6350] <= 1'h0;
      write_enable_data_log_force[6351] <= 1'h0;
      write_enable_data_log_force[6352] <= 1'h0;
      write_enable_data_log_force[6353] <= 1'h0;
      write_enable_data_log_force[6354] <= 1'h0;
      write_enable_data_log_force[6355] <= 1'h0;
      write_enable_data_log_force[6356] <= 1'h0;
      write_enable_data_log_force[6357] <= 1'h0;
      write_enable_data_log_force[6358] <= 1'h0;
      write_enable_data_log_force[6359] <= 1'h0;
      write_enable_data_log_force[6360] <= 1'h0;
      write_enable_data_log_force[6361] <= 1'h0;
      write_enable_data_log_force[6362] <= 1'h0;
      write_enable_data_log_force[6363] <= 1'h0;
      write_enable_data_log_force[6364] <= 1'h0;
      write_enable_data_log_force[6365] <= 1'h0;
      write_enable_data_log_force[6366] <= 1'h0;
      write_enable_data_log_force[6367] <= 1'h0;
      write_enable_data_log_force[6368] <= 1'h0;
      write_enable_data_log_force[6369] <= 1'h0;
      write_enable_data_log_force[6370] <= 1'h0;
      write_enable_data_log_force[6371] <= 1'h0;
      write_enable_data_log_force[6372] <= 1'h0;
      write_enable_data_log_force[6373] <= 1'h0;
      write_enable_data_log_force[6374] <= 1'h0;
      write_enable_data_log_force[6375] <= 1'h0;
      write_enable_data_log_force[6376] <= 1'h0;
      write_enable_data_log_force[6377] <= 1'h0;
      write_enable_data_log_force[6378] <= 1'h0;
      write_enable_data_log_force[6379] <= 1'h0;
      write_enable_data_log_force[6380] <= 1'h0;
      write_enable_data_log_force[6381] <= 1'h0;
      write_enable_data_log_force[6382] <= 1'h0;
      write_enable_data_log_force[6383] <= 1'h0;
      write_enable_data_log_force[6384] <= 1'h0;
      write_enable_data_log_force[6385] <= 1'h0;
      write_enable_data_log_force[6386] <= 1'h0;
      write_enable_data_log_force[6387] <= 1'h0;
      write_enable_data_log_force[6388] <= 1'h0;
      write_enable_data_log_force[6389] <= 1'h0;
      write_enable_data_log_force[6390] <= 1'h0;
      write_enable_data_log_force[6391] <= 1'h0;
      write_enable_data_log_force[6392] <= 1'h0;
      write_enable_data_log_force[6393] <= 1'h0;
      write_enable_data_log_force[6394] <= 1'h0;
      write_enable_data_log_force[6395] <= 1'h0;
      write_enable_data_log_force[6396] <= 1'h0;
      write_enable_data_log_force[6397] <= 1'h0;
      write_enable_data_log_force[6398] <= 1'h0;
      write_enable_data_log_force[6399] <= 1'h0;
      write_enable_data_log_force[6400] <= 1'h0;
      write_enable_data_log_force[6401] <= 1'h0;
      write_enable_data_log_force[6402] <= 1'h0;
      write_enable_data_log_force[6403] <= 1'h0;
      write_enable_data_log_force[6404] <= 1'h0;
      write_enable_data_log_force[6405] <= 1'h0;
      write_enable_data_log_force[6406] <= 1'h0;
      write_enable_data_log_force[6407] <= 1'h0;
      write_enable_data_log_force[6408] <= 1'h0;
      write_enable_data_log_force[6409] <= 1'h0;
      write_enable_data_log_force[6410] <= 1'h0;
      write_enable_data_log_force[6411] <= 1'h0;
      write_enable_data_log_force[6412] <= 1'h0;
      write_enable_data_log_force[6413] <= 1'h0;
      write_enable_data_log_force[6414] <= 1'h0;
      write_enable_data_log_force[6415] <= 1'h0;
      write_enable_data_log_force[6416] <= 1'h0;
      write_enable_data_log_force[6417] <= 1'h0;
      write_enable_data_log_force[6418] <= 1'h0;
      write_enable_data_log_force[6419] <= 1'h0;
      write_enable_data_log_force[6420] <= 1'h0;
      write_enable_data_log_force[6421] <= 1'h0;
      write_enable_data_log_force[6422] <= 1'h0;
      write_enable_data_log_force[6423] <= 1'h0;
      write_enable_data_log_force[6424] <= 1'h0;
      write_enable_data_log_force[6425] <= 1'h0;
      write_enable_data_log_force[6426] <= 1'h0;
      write_enable_data_log_force[6427] <= 1'h0;
      write_enable_data_log_force[6428] <= 1'h0;
      write_enable_data_log_force[6429] <= 1'h0;
      write_enable_data_log_force[6430] <= 1'h0;
      write_enable_data_log_force[6431] <= 1'h0;
      write_enable_data_log_force[6432] <= 1'h0;
      write_enable_data_log_force[6433] <= 1'h0;
      write_enable_data_log_force[6434] <= 1'h0;
      write_enable_data_log_force[6435] <= 1'h0;
      write_enable_data_log_force[6436] <= 1'h0;
      write_enable_data_log_force[6437] <= 1'h0;
      write_enable_data_log_force[6438] <= 1'h0;
      write_enable_data_log_force[6439] <= 1'h0;
      write_enable_data_log_force[6440] <= 1'h0;
      write_enable_data_log_force[6441] <= 1'h0;
      write_enable_data_log_force[6442] <= 1'h0;
      write_enable_data_log_force[6443] <= 1'h0;
      write_enable_data_log_force[6444] <= 1'h0;
      write_enable_data_log_force[6445] <= 1'h0;
      write_enable_data_log_force[6446] <= 1'h0;
      write_enable_data_log_force[6447] <= 1'h0;
      write_enable_data_log_force[6448] <= 1'h0;
      write_enable_data_log_force[6449] <= 1'h0;
      write_enable_data_log_force[6450] <= 1'h0;
      write_enable_data_log_force[6451] <= 1'h0;
      write_enable_data_log_force[6452] <= 1'h0;
      write_enable_data_log_force[6453] <= 1'h0;
      write_enable_data_log_force[6454] <= 1'h0;
      write_enable_data_log_force[6455] <= 1'h0;
      write_enable_data_log_force[6456] <= 1'h0;
      write_enable_data_log_force[6457] <= 1'h0;
      write_enable_data_log_force[6458] <= 1'h0;
      write_enable_data_log_force[6459] <= 1'h0;
      write_enable_data_log_force[6460] <= 1'h0;
      write_enable_data_log_force[6461] <= 1'h0;
      write_enable_data_log_force[6462] <= 1'h0;
      write_enable_data_log_force[6463] <= 1'h0;
      write_enable_data_log_force[6464] <= 1'h0;
      write_enable_data_log_force[6465] <= 1'h0;
      write_enable_data_log_force[6466] <= 1'h0;
      write_enable_data_log_force[6467] <= 1'h0;
      write_enable_data_log_force[6468] <= 1'h0;
      write_enable_data_log_force[6469] <= 1'h0;
      write_enable_data_log_force[6470] <= 1'h0;
      write_enable_data_log_force[6471] <= 1'h0;
      write_enable_data_log_force[6472] <= 1'h0;
      write_enable_data_log_force[6473] <= 1'h0;
      write_enable_data_log_force[6474] <= 1'h0;
      write_enable_data_log_force[6475] <= 1'h0;
      write_enable_data_log_force[6476] <= 1'h0;
      write_enable_data_log_force[6477] <= 1'h0;
      write_enable_data_log_force[6478] <= 1'h0;
      write_enable_data_log_force[6479] <= 1'h0;
      write_enable_data_log_force[6480] <= 1'h0;
      write_enable_data_log_force[6481] <= 1'h0;
      write_enable_data_log_force[6482] <= 1'h0;
      write_enable_data_log_force[6483] <= 1'h0;
      write_enable_data_log_force[6484] <= 1'h0;
      write_enable_data_log_force[6485] <= 1'h0;
      write_enable_data_log_force[6486] <= 1'h0;
      write_enable_data_log_force[6487] <= 1'h0;
      write_enable_data_log_force[6488] <= 1'h0;
      write_enable_data_log_force[6489] <= 1'h0;
      write_enable_data_log_force[6490] <= 1'h0;
      write_enable_data_log_force[6491] <= 1'h0;
      write_enable_data_log_force[6492] <= 1'h0;
      write_enable_data_log_force[6493] <= 1'h0;
      write_enable_data_log_force[6494] <= 1'h0;
      write_enable_data_log_force[6495] <= 1'h0;
      write_enable_data_log_force[6496] <= 1'h0;
      write_enable_data_log_force[6497] <= 1'h0;
      write_enable_data_log_force[6498] <= 1'h0;
      write_enable_data_log_force[6499] <= 1'h0;
      write_enable_data_log_force[6500] <= 1'h0;
      write_enable_data_log_force[6501] <= 1'h0;
      write_enable_data_log_force[6502] <= 1'h0;
      write_enable_data_log_force[6503] <= 1'h0;
      write_enable_data_log_force[6504] <= 1'h0;
      write_enable_data_log_force[6505] <= 1'h0;
      write_enable_data_log_force[6506] <= 1'h0;
      write_enable_data_log_force[6507] <= 1'h0;
      write_enable_data_log_force[6508] <= 1'h0;
      write_enable_data_log_force[6509] <= 1'h0;
      write_enable_data_log_force[6510] <= 1'h0;
      write_enable_data_log_force[6511] <= 1'h0;
      write_enable_data_log_force[6512] <= 1'h0;
      write_enable_data_log_force[6513] <= 1'h0;
      write_enable_data_log_force[6514] <= 1'h0;
      write_enable_data_log_force[6515] <= 1'h0;
      write_enable_data_log_force[6516] <= 1'h0;
      write_enable_data_log_force[6517] <= 1'h0;
      write_enable_data_log_force[6518] <= 1'h0;
      write_enable_data_log_force[6519] <= 1'h0;
      write_enable_data_log_force[6520] <= 1'h0;
      write_enable_data_log_force[6521] <= 1'h0;
      write_enable_data_log_force[6522] <= 1'h0;
      write_enable_data_log_force[6523] <= 1'h0;
      write_enable_data_log_force[6524] <= 1'h0;
      write_enable_data_log_force[6525] <= 1'h0;
      write_enable_data_log_force[6526] <= 1'h0;
      write_enable_data_log_force[6527] <= 1'h0;
      write_enable_data_log_force[6528] <= 1'h0;
      write_enable_data_log_force[6529] <= 1'h0;
      write_enable_data_log_force[6530] <= 1'h0;
      write_enable_data_log_force[6531] <= 1'h0;
      write_enable_data_log_force[6532] <= 1'h0;
      write_enable_data_log_force[6533] <= 1'h0;
      write_enable_data_log_force[6534] <= 1'h0;
      write_enable_data_log_force[6535] <= 1'h0;
      write_enable_data_log_force[6536] <= 1'h0;
      write_enable_data_log_force[6537] <= 1'h0;
      write_enable_data_log_force[6538] <= 1'h0;
      write_enable_data_log_force[6539] <= 1'h0;
      write_enable_data_log_force[6540] <= 1'h0;
      write_enable_data_log_force[6541] <= 1'h0;
      write_enable_data_log_force[6542] <= 1'h0;
      write_enable_data_log_force[6543] <= 1'h0;
      write_enable_data_log_force[6544] <= 1'h0;
      write_enable_data_log_force[6545] <= 1'h0;
      write_enable_data_log_force[6546] <= 1'h0;
      write_enable_data_log_force[6547] <= 1'h0;
      write_enable_data_log_force[6548] <= 1'h0;
      write_enable_data_log_force[6549] <= 1'h0;
      write_enable_data_log_force[6550] <= 1'h0;
      write_enable_data_log_force[6551] <= 1'h0;
      write_enable_data_log_force[6552] <= 1'h0;
      write_enable_data_log_force[6553] <= 1'h0;
      write_enable_data_log_force[6554] <= 1'h0;
      write_enable_data_log_force[6555] <= 1'h0;
      write_enable_data_log_force[6556] <= 1'h0;
      write_enable_data_log_force[6557] <= 1'h0;
      write_enable_data_log_force[6558] <= 1'h0;
      write_enable_data_log_force[6559] <= 1'h0;
      write_enable_data_log_force[6560] <= 1'h0;
      write_enable_data_log_force[6561] <= 1'h0;
      write_enable_data_log_force[6562] <= 1'h0;
      write_enable_data_log_force[6563] <= 1'h0;
      write_enable_data_log_force[6564] <= 1'h0;
      write_enable_data_log_force[6565] <= 1'h0;
      write_enable_data_log_force[6566] <= 1'h0;
      write_enable_data_log_force[6567] <= 1'h0;
      write_enable_data_log_force[6568] <= 1'h0;
      write_enable_data_log_force[6569] <= 1'h0;
      write_enable_data_log_force[6570] <= 1'h0;
      write_enable_data_log_force[6571] <= 1'h0;
      write_enable_data_log_force[6572] <= 1'h0;
      write_enable_data_log_force[6573] <= 1'h0;
      write_enable_data_log_force[6574] <= 1'h0;
      write_enable_data_log_force[6575] <= 1'h0;
      write_enable_data_log_force[6576] <= 1'h0;
      write_enable_data_log_force[6577] <= 1'h0;
      write_enable_data_log_force[6578] <= 1'h0;
      write_enable_data_log_force[6579] <= 1'h0;
      write_enable_data_log_force[6580] <= 1'h0;
      write_enable_data_log_force[6581] <= 1'h0;
      write_enable_data_log_force[6582] <= 1'h0;
      write_enable_data_log_force[6583] <= 1'h0;
      write_enable_data_log_force[6584] <= 1'h0;
      write_enable_data_log_force[6585] <= 1'h0;
      write_enable_data_log_force[6586] <= 1'h0;
      write_enable_data_log_force[6587] <= 1'h0;
      write_enable_data_log_force[6588] <= 1'h0;
      write_enable_data_log_force[6589] <= 1'h0;
      write_enable_data_log_force[6590] <= 1'h0;
      write_enable_data_log_force[6591] <= 1'h0;
      write_enable_data_log_force[6592] <= 1'h0;
      write_enable_data_log_force[6593] <= 1'h0;
      write_enable_data_log_force[6594] <= 1'h0;
      write_enable_data_log_force[6595] <= 1'h0;
      write_enable_data_log_force[6596] <= 1'h0;
      write_enable_data_log_force[6597] <= 1'h0;
      write_enable_data_log_force[6598] <= 1'h0;
      write_enable_data_log_force[6599] <= 1'h0;
      write_enable_data_log_force[6600] <= 1'h0;
      write_enable_data_log_force[6601] <= 1'h0;
      write_enable_data_log_force[6602] <= 1'h0;
      write_enable_data_log_force[6603] <= 1'h0;
      write_enable_data_log_force[6604] <= 1'h0;
      write_enable_data_log_force[6605] <= 1'h0;
      write_enable_data_log_force[6606] <= 1'h0;
      write_enable_data_log_force[6607] <= 1'h0;
      write_enable_data_log_force[6608] <= 1'h0;
      write_enable_data_log_force[6609] <= 1'h0;
      write_enable_data_log_force[6610] <= 1'h0;
      write_enable_data_log_force[6611] <= 1'h0;
      write_enable_data_log_force[6612] <= 1'h0;
      write_enable_data_log_force[6613] <= 1'h0;
      write_enable_data_log_force[6614] <= 1'h0;
      write_enable_data_log_force[6615] <= 1'h0;
      write_enable_data_log_force[6616] <= 1'h0;
      write_enable_data_log_force[6617] <= 1'h0;
      write_enable_data_log_force[6618] <= 1'h0;
      write_enable_data_log_force[6619] <= 1'h0;
      write_enable_data_log_force[6620] <= 1'h0;
      write_enable_data_log_force[6621] <= 1'h0;
      write_enable_data_log_force[6622] <= 1'h0;
      write_enable_data_log_force[6623] <= 1'h0;
      write_enable_data_log_force[6624] <= 1'h0;
      write_enable_data_log_force[6625] <= 1'h0;
      write_enable_data_log_force[6626] <= 1'h0;
      write_enable_data_log_force[6627] <= 1'h0;
      write_enable_data_log_force[6628] <= 1'h0;
      write_enable_data_log_force[6629] <= 1'h0;
      write_enable_data_log_force[6630] <= 1'h0;
      write_enable_data_log_force[6631] <= 1'h0;
      write_enable_data_log_force[6632] <= 1'h0;
      write_enable_data_log_force[6633] <= 1'h0;
      write_enable_data_log_force[6634] <= 1'h0;
      write_enable_data_log_force[6635] <= 1'h0;
      write_enable_data_log_force[6636] <= 1'h0;
      write_enable_data_log_force[6637] <= 1'h0;
      write_enable_data_log_force[6638] <= 1'h0;
      write_enable_data_log_force[6639] <= 1'h0;
      write_enable_data_log_force[6640] <= 1'h0;
      write_enable_data_log_force[6641] <= 1'h0;
      write_enable_data_log_force[6642] <= 1'h0;
      write_enable_data_log_force[6643] <= 1'h0;
      write_enable_data_log_force[6644] <= 1'h0;
      write_enable_data_log_force[6645] <= 1'h0;
      write_enable_data_log_force[6646] <= 1'h0;
      write_enable_data_log_force[6647] <= 1'h0;
      write_enable_data_log_force[6648] <= 1'h0;
      write_enable_data_log_force[6649] <= 1'h0;
      write_enable_data_log_force[6650] <= 1'h0;
      write_enable_data_log_force[6651] <= 1'h0;
      write_enable_data_log_force[6652] <= 1'h0;
      write_enable_data_log_force[6653] <= 1'h0;
      write_enable_data_log_force[6654] <= 1'h0;
      write_enable_data_log_force[6655] <= 1'h0;
      write_enable_data_log_force[6656] <= 1'h0;
      write_enable_data_log_force[6657] <= 1'h0;
      write_enable_data_log_force[6658] <= 1'h0;
      write_enable_data_log_force[6659] <= 1'h0;
      write_enable_data_log_force[6660] <= 1'h0;
      write_enable_data_log_force[6661] <= 1'h0;
      write_enable_data_log_force[6662] <= 1'h0;
      write_enable_data_log_force[6663] <= 1'h0;
      write_enable_data_log_force[6664] <= 1'h0;
      write_enable_data_log_force[6665] <= 1'h0;
      write_enable_data_log_force[6666] <= 1'h0;
      write_enable_data_log_force[6667] <= 1'h0;
      write_enable_data_log_force[6668] <= 1'h0;
      write_enable_data_log_force[6669] <= 1'h0;
      write_enable_data_log_force[6670] <= 1'h0;
      write_enable_data_log_force[6671] <= 1'h0;
      write_enable_data_log_force[6672] <= 1'h0;
      write_enable_data_log_force[6673] <= 1'h0;
      write_enable_data_log_force[6674] <= 1'h0;
      write_enable_data_log_force[6675] <= 1'h0;
      write_enable_data_log_force[6676] <= 1'h0;
      write_enable_data_log_force[6677] <= 1'h0;
      write_enable_data_log_force[6678] <= 1'h0;
      write_enable_data_log_force[6679] <= 1'h0;
      write_enable_data_log_force[6680] <= 1'h0;
      write_enable_data_log_force[6681] <= 1'h0;
      write_enable_data_log_force[6682] <= 1'h0;
      write_enable_data_log_force[6683] <= 1'h0;
      write_enable_data_log_force[6684] <= 1'h0;
      write_enable_data_log_force[6685] <= 1'h0;
      write_enable_data_log_force[6686] <= 1'h0;
      write_enable_data_log_force[6687] <= 1'h0;
      write_enable_data_log_force[6688] <= 1'h0;
      write_enable_data_log_force[6689] <= 1'h0;
      write_enable_data_log_force[6690] <= 1'h0;
      write_enable_data_log_force[6691] <= 1'h0;
      write_enable_data_log_force[6692] <= 1'h0;
      write_enable_data_log_force[6693] <= 1'h0;
      write_enable_data_log_force[6694] <= 1'h0;
      write_enable_data_log_force[6695] <= 1'h0;
      write_enable_data_log_force[6696] <= 1'h0;
      write_enable_data_log_force[6697] <= 1'h0;
      write_enable_data_log_force[6698] <= 1'h0;
      write_enable_data_log_force[6699] <= 1'h0;
      write_enable_data_log_force[6700] <= 1'h0;
      write_enable_data_log_force[6701] <= 1'h0;
      write_enable_data_log_force[6702] <= 1'h0;
      write_enable_data_log_force[6703] <= 1'h0;
      write_enable_data_log_force[6704] <= 1'h0;
      write_enable_data_log_force[6705] <= 1'h0;
      write_enable_data_log_force[6706] <= 1'h0;
      write_enable_data_log_force[6707] <= 1'h0;
      write_enable_data_log_force[6708] <= 1'h0;
      write_enable_data_log_force[6709] <= 1'h0;
      write_enable_data_log_force[6710] <= 1'h0;
      write_enable_data_log_force[6711] <= 1'h0;
      write_enable_data_log_force[6712] <= 1'h0;
      write_enable_data_log_force[6713] <= 1'h0;
      write_enable_data_log_force[6714] <= 1'h0;
      write_enable_data_log_force[6715] <= 1'h0;
      write_enable_data_log_force[6716] <= 1'h0;
      write_enable_data_log_force[6717] <= 1'h0;
      write_enable_data_log_force[6718] <= 1'h0;
      write_enable_data_log_force[6719] <= 1'h0;
      write_enable_data_log_force[6720] <= 1'h0;
      write_enable_data_log_force[6721] <= 1'h0;
      write_enable_data_log_force[6722] <= 1'h0;
      write_enable_data_log_force[6723] <= 1'h0;
      write_enable_data_log_force[6724] <= 1'h0;
      write_enable_data_log_force[6725] <= 1'h0;
      write_enable_data_log_force[6726] <= 1'h0;
      write_enable_data_log_force[6727] <= 1'h0;
      write_enable_data_log_force[6728] <= 1'h0;
      write_enable_data_log_force[6729] <= 1'h0;
      write_enable_data_log_force[6730] <= 1'h0;
      write_enable_data_log_force[6731] <= 1'h0;
      write_enable_data_log_force[6732] <= 1'h0;
      write_enable_data_log_force[6733] <= 1'h0;
      write_enable_data_log_force[6734] <= 1'h0;
      write_enable_data_log_force[6735] <= 1'h0;
      write_enable_data_log_force[6736] <= 1'h0;
      write_enable_data_log_force[6737] <= 1'h0;
      write_enable_data_log_force[6738] <= 1'h0;
      write_enable_data_log_force[6739] <= 1'h0;
      write_enable_data_log_force[6740] <= 1'h0;
      write_enable_data_log_force[6741] <= 1'h0;
      write_enable_data_log_force[6742] <= 1'h0;
      write_enable_data_log_force[6743] <= 1'h0;
      write_enable_data_log_force[6744] <= 1'h0;
      write_enable_data_log_force[6745] <= 1'h0;
      write_enable_data_log_force[6746] <= 1'h0;
      write_enable_data_log_force[6747] <= 1'h0;
      write_enable_data_log_force[6748] <= 1'h0;
      write_enable_data_log_force[6749] <= 1'h0;
      write_enable_data_log_force[6750] <= 1'h0;
      write_enable_data_log_force[6751] <= 1'h0;
      write_enable_data_log_force[6752] <= 1'h0;
      write_enable_data_log_force[6753] <= 1'h0;
      write_enable_data_log_force[6754] <= 1'h0;
      write_enable_data_log_force[6755] <= 1'h0;
      write_enable_data_log_force[6756] <= 1'h0;
      write_enable_data_log_force[6757] <= 1'h0;
      write_enable_data_log_force[6758] <= 1'h0;
      write_enable_data_log_force[6759] <= 1'h0;
      write_enable_data_log_force[6760] <= 1'h0;
      write_enable_data_log_force[6761] <= 1'h0;
      write_enable_data_log_force[6762] <= 1'h0;
      write_enable_data_log_force[6763] <= 1'h0;
      write_enable_data_log_force[6764] <= 1'h0;
      write_enable_data_log_force[6765] <= 1'h0;
      write_enable_data_log_force[6766] <= 1'h0;
      write_enable_data_log_force[6767] <= 1'h0;
      write_enable_data_log_force[6768] <= 1'h0;
      write_enable_data_log_force[6769] <= 1'h0;
      write_enable_data_log_force[6770] <= 1'h0;
      write_enable_data_log_force[6771] <= 1'h0;
      write_enable_data_log_force[6772] <= 1'h0;
      write_enable_data_log_force[6773] <= 1'h0;
      write_enable_data_log_force[6774] <= 1'h0;
      write_enable_data_log_force[6775] <= 1'h0;
      write_enable_data_log_force[6776] <= 1'h0;
      write_enable_data_log_force[6777] <= 1'h0;
      write_enable_data_log_force[6778] <= 1'h0;
      write_enable_data_log_force[6779] <= 1'h0;
      write_enable_data_log_force[6780] <= 1'h0;
      write_enable_data_log_force[6781] <= 1'h0;
      write_enable_data_log_force[6782] <= 1'h0;
      write_enable_data_log_force[6783] <= 1'h0;
      write_enable_data_log_force[6784] <= 1'h0;
      write_enable_data_log_force[6785] <= 1'h0;
      write_enable_data_log_force[6786] <= 1'h0;
      write_enable_data_log_force[6787] <= 1'h0;
      write_enable_data_log_force[6788] <= 1'h0;
      write_enable_data_log_force[6789] <= 1'h0;
      write_enable_data_log_force[6790] <= 1'h0;
      write_enable_data_log_force[6791] <= 1'h0;
      write_enable_data_log_force[6792] <= 1'h0;
      write_enable_data_log_force[6793] <= 1'h0;
      write_enable_data_log_force[6794] <= 1'h0;
      write_enable_data_log_force[6795] <= 1'h0;
      write_enable_data_log_force[6796] <= 1'h0;
      write_enable_data_log_force[6797] <= 1'h0;
      write_enable_data_log_force[6798] <= 1'h0;
      write_enable_data_log_force[6799] <= 1'h0;
      write_enable_data_log_force[6800] <= 1'h0;
      write_enable_data_log_force[6801] <= 1'h0;
      write_enable_data_log_force[6802] <= 1'h0;
      write_enable_data_log_force[6803] <= 1'h0;
      write_enable_data_log_force[6804] <= 1'h0;
      write_enable_data_log_force[6805] <= 1'h0;
      write_enable_data_log_force[6806] <= 1'h0;
      write_enable_data_log_force[6807] <= 1'h0;
      write_enable_data_log_force[6808] <= 1'h0;
      write_enable_data_log_force[6809] <= 1'h0;
      write_enable_data_log_force[6810] <= 1'h0;
      write_enable_data_log_force[6811] <= 1'h0;
      write_enable_data_log_force[6812] <= 1'h0;
      write_enable_data_log_force[6813] <= 1'h0;
      write_enable_data_log_force[6814] <= 1'h0;
      write_enable_data_log_force[6815] <= 1'h0;
      write_enable_data_log_force[6816] <= 1'h0;
      write_enable_data_log_force[6817] <= 1'h0;
      write_enable_data_log_force[6818] <= 1'h0;
      write_enable_data_log_force[6819] <= 1'h0;
      write_enable_data_log_force[6820] <= 1'h0;
      write_enable_data_log_force[6821] <= 1'h0;
      write_enable_data_log_force[6822] <= 1'h0;
      write_enable_data_log_force[6823] <= 1'h0;
      write_enable_data_log_force[6824] <= 1'h0;
      write_enable_data_log_force[6825] <= 1'h0;
      write_enable_data_log_force[6826] <= 1'h0;
      write_enable_data_log_force[6827] <= 1'h0;
      write_enable_data_log_force[6828] <= 1'h0;
      write_enable_data_log_force[6829] <= 1'h0;
      write_enable_data_log_force[6830] <= 1'h0;
      write_enable_data_log_force[6831] <= 1'h0;
      write_enable_data_log_force[6832] <= 1'h0;
      write_enable_data_log_force[6833] <= 1'h0;
      write_enable_data_log_force[6834] <= 1'h0;
      write_enable_data_log_force[6835] <= 1'h0;
      write_enable_data_log_force[6836] <= 1'h0;
      write_enable_data_log_force[6837] <= 1'h0;
      write_enable_data_log_force[6838] <= 1'h0;
      write_enable_data_log_force[6839] <= 1'h0;
      write_enable_data_log_force[6840] <= 1'h0;
      write_enable_data_log_force[6841] <= 1'h0;
      write_enable_data_log_force[6842] <= 1'h0;
      write_enable_data_log_force[6843] <= 1'h0;
      write_enable_data_log_force[6844] <= 1'h0;
      write_enable_data_log_force[6845] <= 1'h0;
      write_enable_data_log_force[6846] <= 1'h0;
      write_enable_data_log_force[6847] <= 1'h0;
      write_enable_data_log_force[6848] <= 1'h0;
      write_enable_data_log_force[6849] <= 1'h0;
      write_enable_data_log_force[6850] <= 1'h0;
      write_enable_data_log_force[6851] <= 1'h0;
      write_enable_data_log_force[6852] <= 1'h0;
      write_enable_data_log_force[6853] <= 1'h0;
      write_enable_data_log_force[6854] <= 1'h0;
      write_enable_data_log_force[6855] <= 1'h0;
      write_enable_data_log_force[6856] <= 1'h0;
      write_enable_data_log_force[6857] <= 1'h0;
      write_enable_data_log_force[6858] <= 1'h0;
      write_enable_data_log_force[6859] <= 1'h0;
      write_enable_data_log_force[6860] <= 1'h0;
      write_enable_data_log_force[6861] <= 1'h0;
      write_enable_data_log_force[6862] <= 1'h0;
      write_enable_data_log_force[6863] <= 1'h0;
      write_enable_data_log_force[6864] <= 1'h0;
      write_enable_data_log_force[6865] <= 1'h0;
      write_enable_data_log_force[6866] <= 1'h0;
      write_enable_data_log_force[6867] <= 1'h0;
      write_enable_data_log_force[6868] <= 1'h0;
      write_enable_data_log_force[6869] <= 1'h0;
      write_enable_data_log_force[6870] <= 1'h0;
      write_enable_data_log_force[6871] <= 1'h0;
      write_enable_data_log_force[6872] <= 1'h0;
      write_enable_data_log_force[6873] <= 1'h0;
      write_enable_data_log_force[6874] <= 1'h0;
      write_enable_data_log_force[6875] <= 1'h0;
      write_enable_data_log_force[6876] <= 1'h0;
      write_enable_data_log_force[6877] <= 1'h0;
      write_enable_data_log_force[6878] <= 1'h0;
      write_enable_data_log_force[6879] <= 1'h0;
      write_enable_data_log_force[6880] <= 1'h0;
      write_enable_data_log_force[6881] <= 1'h0;
      write_enable_data_log_force[6882] <= 1'h0;
      write_enable_data_log_force[6883] <= 1'h0;
      write_enable_data_log_force[6884] <= 1'h0;
      write_enable_data_log_force[6885] <= 1'h0;
      write_enable_data_log_force[6886] <= 1'h0;
      write_enable_data_log_force[6887] <= 1'h0;
      write_enable_data_log_force[6888] <= 1'h0;
      write_enable_data_log_force[6889] <= 1'h0;
      write_enable_data_log_force[6890] <= 1'h0;
      write_enable_data_log_force[6891] <= 1'h0;
      write_enable_data_log_force[6892] <= 1'h0;
      write_enable_data_log_force[6893] <= 1'h0;
      write_enable_data_log_force[6894] <= 1'h0;
      write_enable_data_log_force[6895] <= 1'h0;
      write_enable_data_log_force[6896] <= 1'h0;
      write_enable_data_log_force[6897] <= 1'h0;
      write_enable_data_log_force[6898] <= 1'h0;
      write_enable_data_log_force[6899] <= 1'h0;
      write_enable_data_log_force[6900] <= 1'h0;
      write_enable_data_log_force[6901] <= 1'h0;
      write_enable_data_log_force[6902] <= 1'h0;
      write_enable_data_log_force[6903] <= 1'h0;
      write_enable_data_log_force[6904] <= 1'h0;
      write_enable_data_log_force[6905] <= 1'h0;
      write_enable_data_log_force[6906] <= 1'h0;
      write_enable_data_log_force[6907] <= 1'h0;
      write_enable_data_log_force[6908] <= 1'h0;
      write_enable_data_log_force[6909] <= 1'h0;
      write_enable_data_log_force[6910] <= 1'h0;
      write_enable_data_log_force[6911] <= 1'h0;
      write_enable_data_log_force[6912] <= 1'h0;
      write_enable_data_log_force[6913] <= 1'h0;
      write_enable_data_log_force[6914] <= 1'h0;
      write_enable_data_log_force[6915] <= 1'h0;
      write_enable_data_log_force[6916] <= 1'h0;
      write_enable_data_log_force[6917] <= 1'h0;
      write_enable_data_log_force[6918] <= 1'h0;
      write_enable_data_log_force[6919] <= 1'h0;
      write_enable_data_log_force[6920] <= 1'h0;
      write_enable_data_log_force[6921] <= 1'h0;
      write_enable_data_log_force[6922] <= 1'h0;
      write_enable_data_log_force[6923] <= 1'h0;
      write_enable_data_log_force[6924] <= 1'h0;
      write_enable_data_log_force[6925] <= 1'h0;
      write_enable_data_log_force[6926] <= 1'h0;
      write_enable_data_log_force[6927] <= 1'h0;
      write_enable_data_log_force[6928] <= 1'h0;
      write_enable_data_log_force[6929] <= 1'h0;
      write_enable_data_log_force[6930] <= 1'h0;
      write_enable_data_log_force[6931] <= 1'h0;
      write_enable_data_log_force[6932] <= 1'h0;
      write_enable_data_log_force[6933] <= 1'h0;
      write_enable_data_log_force[6934] <= 1'h0;
      write_enable_data_log_force[6935] <= 1'h0;
      write_enable_data_log_force[6936] <= 1'h0;
      write_enable_data_log_force[6937] <= 1'h0;
      write_enable_data_log_force[6938] <= 1'h0;
      write_enable_data_log_force[6939] <= 1'h0;
      write_enable_data_log_force[6940] <= 1'h0;
      write_enable_data_log_force[6941] <= 1'h0;
      write_enable_data_log_force[6942] <= 1'h0;
      write_enable_data_log_force[6943] <= 1'h0;
      write_enable_data_log_force[6944] <= 1'h0;
      write_enable_data_log_force[6945] <= 1'h0;
      write_enable_data_log_force[6946] <= 1'h0;
      write_enable_data_log_force[6947] <= 1'h0;
      write_enable_data_log_force[6948] <= 1'h0;
      write_enable_data_log_force[6949] <= 1'h0;
      write_enable_data_log_force[6950] <= 1'h0;
      write_enable_data_log_force[6951] <= 1'h0;
      write_enable_data_log_force[6952] <= 1'h0;
      write_enable_data_log_force[6953] <= 1'h0;
      write_enable_data_log_force[6954] <= 1'h0;
      write_enable_data_log_force[6955] <= 1'h0;
      write_enable_data_log_force[6956] <= 1'h0;
      write_enable_data_log_force[6957] <= 1'h0;
      write_enable_data_log_force[6958] <= 1'h0;
      write_enable_data_log_force[6959] <= 1'h0;
      write_enable_data_log_force[6960] <= 1'h0;
      write_enable_data_log_force[6961] <= 1'h0;
      write_enable_data_log_force[6962] <= 1'h0;
      write_enable_data_log_force[6963] <= 1'h0;
      write_enable_data_log_force[6964] <= 1'h0;
      write_enable_data_log_force[6965] <= 1'h0;
      write_enable_data_log_force[6966] <= 1'h0;
      write_enable_data_log_force[6967] <= 1'h0;
      write_enable_data_log_force[6968] <= 1'h0;
      write_enable_data_log_force[6969] <= 1'h0;
      write_enable_data_log_force[6970] <= 1'h0;
      write_enable_data_log_force[6971] <= 1'h0;
      write_enable_data_log_force[6972] <= 1'h0;
      write_enable_data_log_force[6973] <= 1'h0;
      write_enable_data_log_force[6974] <= 1'h0;
      write_enable_data_log_force[6975] <= 1'h0;
      write_enable_data_log_force[6976] <= 1'h0;
      write_enable_data_log_force[6977] <= 1'h0;
      write_enable_data_log_force[6978] <= 1'h0;
      write_enable_data_log_force[6979] <= 1'h0;
      write_enable_data_log_force[6980] <= 1'h0;
      write_enable_data_log_force[6981] <= 1'h0;
      write_enable_data_log_force[6982] <= 1'h0;
      write_enable_data_log_force[6983] <= 1'h0;
      write_enable_data_log_force[6984] <= 1'h0;
      write_enable_data_log_force[6985] <= 1'h0;
      write_enable_data_log_force[6986] <= 1'h0;
      write_enable_data_log_force[6987] <= 1'h0;
      write_enable_data_log_force[6988] <= 1'h0;
      write_enable_data_log_force[6989] <= 1'h0;
      write_enable_data_log_force[6990] <= 1'h0;
      write_enable_data_log_force[6991] <= 1'h0;
      write_enable_data_log_force[6992] <= 1'h0;
      write_enable_data_log_force[6993] <= 1'h0;
      write_enable_data_log_force[6994] <= 1'h0;
      write_enable_data_log_force[6995] <= 1'h0;
      write_enable_data_log_force[6996] <= 1'h0;
      write_enable_data_log_force[6997] <= 1'h0;
      write_enable_data_log_force[6998] <= 1'h0;
      write_enable_data_log_force[6999] <= 1'h0;
      write_enable_data_log_force[7000] <= 1'h0;
      write_enable_data_log_force[7001] <= 1'h0;
      write_enable_data_log_force[7002] <= 1'h0;
      write_enable_data_log_force[7003] <= 1'h0;
      write_enable_data_log_force[7004] <= 1'h0;
      write_enable_data_log_force[7005] <= 1'h0;
      write_enable_data_log_force[7006] <= 1'h0;
      write_enable_data_log_force[7007] <= 1'h0;
      write_enable_data_log_force[7008] <= 1'h0;
      write_enable_data_log_force[7009] <= 1'h0;
      write_enable_data_log_force[7010] <= 1'h0;
      write_enable_data_log_force[7011] <= 1'h0;
      write_enable_data_log_force[7012] <= 1'h0;
      write_enable_data_log_force[7013] <= 1'h0;
      write_enable_data_log_force[7014] <= 1'h0;
      write_enable_data_log_force[7015] <= 1'h0;
      write_enable_data_log_force[7016] <= 1'h0;
      write_enable_data_log_force[7017] <= 1'h0;
      write_enable_data_log_force[7018] <= 1'h0;
      write_enable_data_log_force[7019] <= 1'h0;
      write_enable_data_log_force[7020] <= 1'h0;
      write_enable_data_log_force[7021] <= 1'h0;
      write_enable_data_log_force[7022] <= 1'h0;
      write_enable_data_log_force[7023] <= 1'h0;
      write_enable_data_log_force[7024] <= 1'h0;
      write_enable_data_log_force[7025] <= 1'h0;
      write_enable_data_log_force[7026] <= 1'h0;
      write_enable_data_log_force[7027] <= 1'h0;
      write_enable_data_log_force[7028] <= 1'h0;
      write_enable_data_log_force[7029] <= 1'h0;
      write_enable_data_log_force[7030] <= 1'h0;
      write_enable_data_log_force[7031] <= 1'h0;
      write_enable_data_log_force[7032] <= 1'h0;
      write_enable_data_log_force[7033] <= 1'h0;
      write_enable_data_log_force[7034] <= 1'h0;
      write_enable_data_log_force[7035] <= 1'h0;
      write_enable_data_log_force[7036] <= 1'h0;
      write_enable_data_log_force[7037] <= 1'h0;
      write_enable_data_log_force[7038] <= 1'h0;
      write_enable_data_log_force[7039] <= 1'h0;
      write_enable_data_log_force[7040] <= 1'h0;
      write_enable_data_log_force[7041] <= 1'h0;
      write_enable_data_log_force[7042] <= 1'h0;
      write_enable_data_log_force[7043] <= 1'h0;
      write_enable_data_log_force[7044] <= 1'h0;
      write_enable_data_log_force[7045] <= 1'h0;
      write_enable_data_log_force[7046] <= 1'h0;
      write_enable_data_log_force[7047] <= 1'h0;
      write_enable_data_log_force[7048] <= 1'h0;
      write_enable_data_log_force[7049] <= 1'h0;
      write_enable_data_log_force[7050] <= 1'h0;
      write_enable_data_log_force[7051] <= 1'h0;
      write_enable_data_log_force[7052] <= 1'h0;
      write_enable_data_log_force[7053] <= 1'h0;
      write_enable_data_log_force[7054] <= 1'h0;
      write_enable_data_log_force[7055] <= 1'h0;
      write_enable_data_log_force[7056] <= 1'h0;
      write_enable_data_log_force[7057] <= 1'h0;
      write_enable_data_log_force[7058] <= 1'h0;
      write_enable_data_log_force[7059] <= 1'h0;
      write_enable_data_log_force[7060] <= 1'h0;
      write_enable_data_log_force[7061] <= 1'h0;
      write_enable_data_log_force[7062] <= 1'h0;
      write_enable_data_log_force[7063] <= 1'h0;
      write_enable_data_log_force[7064] <= 1'h0;
      write_enable_data_log_force[7065] <= 1'h0;
      write_enable_data_log_force[7066] <= 1'h0;
      write_enable_data_log_force[7067] <= 1'h0;
      write_enable_data_log_force[7068] <= 1'h0;
      write_enable_data_log_force[7069] <= 1'h0;
      write_enable_data_log_force[7070] <= 1'h0;
      write_enable_data_log_force[7071] <= 1'h0;
      write_enable_data_log_force[7072] <= 1'h0;
      write_enable_data_log_force[7073] <= 1'h0;
      write_enable_data_log_force[7074] <= 1'h0;
      write_enable_data_log_force[7075] <= 1'h0;
      write_enable_data_log_force[7076] <= 1'h0;
      write_enable_data_log_force[7077] <= 1'h0;
      write_enable_data_log_force[7078] <= 1'h0;
      write_enable_data_log_force[7079] <= 1'h0;
      write_enable_data_log_force[7080] <= 1'h0;
      write_enable_data_log_force[7081] <= 1'h0;
      write_enable_data_log_force[7082] <= 1'h0;
      write_enable_data_log_force[7083] <= 1'h0;
      write_enable_data_log_force[7084] <= 1'h0;
      write_enable_data_log_force[7085] <= 1'h0;
      write_enable_data_log_force[7086] <= 1'h0;
      write_enable_data_log_force[7087] <= 1'h0;
      write_enable_data_log_force[7088] <= 1'h0;
      write_enable_data_log_force[7089] <= 1'h0;
      write_enable_data_log_force[7090] <= 1'h0;
      write_enable_data_log_force[7091] <= 1'h0;
      write_enable_data_log_force[7092] <= 1'h0;
      write_enable_data_log_force[7093] <= 1'h0;
      write_enable_data_log_force[7094] <= 1'h0;
      write_enable_data_log_force[7095] <= 1'h0;
      write_enable_data_log_force[7096] <= 1'h0;
      write_enable_data_log_force[7097] <= 1'h0;
      write_enable_data_log_force[7098] <= 1'h0;
      write_enable_data_log_force[7099] <= 1'h0;
      write_enable_data_log_force[7100] <= 1'h0;
      write_enable_data_log_force[7101] <= 1'h0;
      write_enable_data_log_force[7102] <= 1'h0;
      write_enable_data_log_force[7103] <= 1'h0;
      write_enable_data_log_force[7104] <= 1'h0;
      write_enable_data_log_force[7105] <= 1'h0;
      write_enable_data_log_force[7106] <= 1'h0;
      write_enable_data_log_force[7107] <= 1'h0;
      write_enable_data_log_force[7108] <= 1'h0;
      write_enable_data_log_force[7109] <= 1'h0;
      write_enable_data_log_force[7110] <= 1'h0;
      write_enable_data_log_force[7111] <= 1'h0;
      write_enable_data_log_force[7112] <= 1'h0;
      write_enable_data_log_force[7113] <= 1'h0;
      write_enable_data_log_force[7114] <= 1'h0;
      write_enable_data_log_force[7115] <= 1'h0;
      write_enable_data_log_force[7116] <= 1'h0;
      write_enable_data_log_force[7117] <= 1'h0;
      write_enable_data_log_force[7118] <= 1'h0;
      write_enable_data_log_force[7119] <= 1'h0;
      write_enable_data_log_force[7120] <= 1'h0;
      write_enable_data_log_force[7121] <= 1'h0;
      write_enable_data_log_force[7122] <= 1'h0;
      write_enable_data_log_force[7123] <= 1'h0;
      write_enable_data_log_force[7124] <= 1'h0;
      write_enable_data_log_force[7125] <= 1'h0;
      write_enable_data_log_force[7126] <= 1'h0;
      write_enable_data_log_force[7127] <= 1'h0;
      write_enable_data_log_force[7128] <= 1'h0;
      write_enable_data_log_force[7129] <= 1'h0;
      write_enable_data_log_force[7130] <= 1'h0;
      write_enable_data_log_force[7131] <= 1'h0;
      write_enable_data_log_force[7132] <= 1'h0;
      write_enable_data_log_force[7133] <= 1'h0;
      write_enable_data_log_force[7134] <= 1'h0;
      write_enable_data_log_force[7135] <= 1'h0;
      write_enable_data_log_force[7136] <= 1'h0;
      write_enable_data_log_force[7137] <= 1'h0;
      write_enable_data_log_force[7138] <= 1'h0;
      write_enable_data_log_force[7139] <= 1'h0;
      write_enable_data_log_force[7140] <= 1'h0;
      write_enable_data_log_force[7141] <= 1'h0;
      write_enable_data_log_force[7142] <= 1'h0;
      write_enable_data_log_force[7143] <= 1'h0;
      write_enable_data_log_force[7144] <= 1'h0;
      write_enable_data_log_force[7145] <= 1'h0;
      write_enable_data_log_force[7146] <= 1'h0;
      write_enable_data_log_force[7147] <= 1'h0;
      write_enable_data_log_force[7148] <= 1'h0;
      write_enable_data_log_force[7149] <= 1'h0;
      write_enable_data_log_force[7150] <= 1'h0;
      write_enable_data_log_force[7151] <= 1'h0;
      write_enable_data_log_force[7152] <= 1'h0;
      write_enable_data_log_force[7153] <= 1'h0;
      write_enable_data_log_force[7154] <= 1'h0;
      write_enable_data_log_force[7155] <= 1'h0;
      write_enable_data_log_force[7156] <= 1'h0;
      write_enable_data_log_force[7157] <= 1'h0;
      write_enable_data_log_force[7158] <= 1'h0;
      write_enable_data_log_force[7159] <= 1'h0;
      write_enable_data_log_force[7160] <= 1'h0;
      write_enable_data_log_force[7161] <= 1'h0;
      write_enable_data_log_force[7162] <= 1'h0;
      write_enable_data_log_force[7163] <= 1'h0;
      write_enable_data_log_force[7164] <= 1'h0;
      write_enable_data_log_force[7165] <= 1'h0;
      write_enable_data_log_force[7166] <= 1'h0;
      write_enable_data_log_force[7167] <= 1'h0;
      write_enable_data_log_force[7168] <= 1'h0;
      write_enable_data_log_force[7169] <= 1'h0;
      write_enable_data_log_force[7170] <= 1'h0;
      write_enable_data_log_force[7171] <= 1'h0;
      write_enable_data_log_force[7172] <= 1'h0;
      write_enable_data_log_force[7173] <= 1'h0;
      write_enable_data_log_force[7174] <= 1'h0;
      write_enable_data_log_force[7175] <= 1'h0;
      write_enable_data_log_force[7176] <= 1'h0;
      write_enable_data_log_force[7177] <= 1'h0;
      write_enable_data_log_force[7178] <= 1'h0;
      write_enable_data_log_force[7179] <= 1'h0;
      write_enable_data_log_force[7180] <= 1'h0;
      write_enable_data_log_force[7181] <= 1'h0;
      write_enable_data_log_force[7182] <= 1'h0;
      write_enable_data_log_force[7183] <= 1'h0;
      write_enable_data_log_force[7184] <= 1'h0;
      write_enable_data_log_force[7185] <= 1'h0;
      write_enable_data_log_force[7186] <= 1'h0;
      write_enable_data_log_force[7187] <= 1'h0;
      write_enable_data_log_force[7188] <= 1'h0;
      write_enable_data_log_force[7189] <= 1'h0;
      write_enable_data_log_force[7190] <= 1'h0;
      write_enable_data_log_force[7191] <= 1'h0;
      write_enable_data_log_force[7192] <= 1'h0;
      write_enable_data_log_force[7193] <= 1'h0;
      write_enable_data_log_force[7194] <= 1'h0;
      write_enable_data_log_force[7195] <= 1'h0;
      write_enable_data_log_force[7196] <= 1'h0;
      write_enable_data_log_force[7197] <= 1'h0;
      write_enable_data_log_force[7198] <= 1'h0;
      write_enable_data_log_force[7199] <= 1'h0;
      write_enable_data_log_force[7200] <= 1'h0;
      write_enable_data_log_force[7201] <= 1'h0;
      write_enable_data_log_force[7202] <= 1'h0;
      write_enable_data_log_force[7203] <= 1'h0;
      write_enable_data_log_force[7204] <= 1'h0;
      write_enable_data_log_force[7205] <= 1'h0;
      write_enable_data_log_force[7206] <= 1'h0;
      write_enable_data_log_force[7207] <= 1'h0;
      write_enable_data_log_force[7208] <= 1'h0;
      write_enable_data_log_force[7209] <= 1'h0;
      write_enable_data_log_force[7210] <= 1'h0;
      write_enable_data_log_force[7211] <= 1'h0;
      write_enable_data_log_force[7212] <= 1'h0;
      write_enable_data_log_force[7213] <= 1'h0;
      write_enable_data_log_force[7214] <= 1'h0;
      write_enable_data_log_force[7215] <= 1'h0;
      write_enable_data_log_force[7216] <= 1'h0;
      write_enable_data_log_force[7217] <= 1'h0;
      write_enable_data_log_force[7218] <= 1'h0;
      write_enable_data_log_force[7219] <= 1'h0;
      write_enable_data_log_force[7220] <= 1'h0;
      write_enable_data_log_force[7221] <= 1'h0;
      write_enable_data_log_force[7222] <= 1'h0;
      write_enable_data_log_force[7223] <= 1'h0;
      write_enable_data_log_force[7224] <= 1'h0;
      write_enable_data_log_force[7225] <= 1'h0;
      write_enable_data_log_force[7226] <= 1'h0;
      write_enable_data_log_force[7227] <= 1'h0;
      write_enable_data_log_force[7228] <= 1'h0;
      write_enable_data_log_force[7229] <= 1'h0;
      write_enable_data_log_force[7230] <= 1'h0;
      write_enable_data_log_force[7231] <= 1'h0;
      write_enable_data_log_force[7232] <= 1'h0;
      write_enable_data_log_force[7233] <= 1'h0;
      write_enable_data_log_force[7234] <= 1'h0;
      write_enable_data_log_force[7235] <= 1'h0;
      write_enable_data_log_force[7236] <= 1'h0;
      write_enable_data_log_force[7237] <= 1'h0;
      write_enable_data_log_force[7238] <= 1'h0;
      write_enable_data_log_force[7239] <= 1'h0;
      write_enable_data_log_force[7240] <= 1'h0;
      write_enable_data_log_force[7241] <= 1'h0;
      write_enable_data_log_force[7242] <= 1'h0;
      write_enable_data_log_force[7243] <= 1'h0;
      write_enable_data_log_force[7244] <= 1'h0;
      write_enable_data_log_force[7245] <= 1'h0;
      write_enable_data_log_force[7246] <= 1'h0;
      write_enable_data_log_force[7247] <= 1'h0;
      write_enable_data_log_force[7248] <= 1'h0;
      write_enable_data_log_force[7249] <= 1'h0;
      write_enable_data_log_force[7250] <= 1'h0;
      write_enable_data_log_force[7251] <= 1'h0;
      write_enable_data_log_force[7252] <= 1'h0;
      write_enable_data_log_force[7253] <= 1'h0;
      write_enable_data_log_force[7254] <= 1'h0;
      write_enable_data_log_force[7255] <= 1'h0;
      write_enable_data_log_force[7256] <= 1'h0;
      write_enable_data_log_force[7257] <= 1'h0;
      write_enable_data_log_force[7258] <= 1'h0;
      write_enable_data_log_force[7259] <= 1'h0;
      write_enable_data_log_force[7260] <= 1'h0;
      write_enable_data_log_force[7261] <= 1'h0;
      write_enable_data_log_force[7262] <= 1'h0;
      write_enable_data_log_force[7263] <= 1'h0;
      write_enable_data_log_force[7264] <= 1'h0;
      write_enable_data_log_force[7265] <= 1'h0;
      write_enable_data_log_force[7266] <= 1'h0;
      write_enable_data_log_force[7267] <= 1'h0;
      write_enable_data_log_force[7268] <= 1'h0;
      write_enable_data_log_force[7269] <= 1'h0;
      write_enable_data_log_force[7270] <= 1'h0;
      write_enable_data_log_force[7271] <= 1'h0;
      write_enable_data_log_force[7272] <= 1'h0;
      write_enable_data_log_force[7273] <= 1'h0;
      write_enable_data_log_force[7274] <= 1'h0;
      write_enable_data_log_force[7275] <= 1'h0;
      write_enable_data_log_force[7276] <= 1'h0;
      write_enable_data_log_force[7277] <= 1'h0;
      write_enable_data_log_force[7278] <= 1'h0;
      write_enable_data_log_force[7279] <= 1'h0;
      write_enable_data_log_force[7280] <= 1'h0;
      write_enable_data_log_force[7281] <= 1'h0;
      write_enable_data_log_force[7282] <= 1'h0;
      write_enable_data_log_force[7283] <= 1'h0;
      write_enable_data_log_force[7284] <= 1'h0;
      write_enable_data_log_force[7285] <= 1'h0;
      write_enable_data_log_force[7286] <= 1'h0;
      write_enable_data_log_force[7287] <= 1'h0;
      write_enable_data_log_force[7288] <= 1'h0;
      write_enable_data_log_force[7289] <= 1'h0;
      write_enable_data_log_force[7290] <= 1'h0;
      write_enable_data_log_force[7291] <= 1'h0;
      write_enable_data_log_force[7292] <= 1'h0;
      write_enable_data_log_force[7293] <= 1'h0;
      write_enable_data_log_force[7294] <= 1'h0;
      write_enable_data_log_force[7295] <= 1'h0;
      write_enable_data_log_force[7296] <= 1'h0;
      write_enable_data_log_force[7297] <= 1'h0;
      write_enable_data_log_force[7298] <= 1'h0;
      write_enable_data_log_force[7299] <= 1'h0;
      write_enable_data_log_force[7300] <= 1'h0;
      write_enable_data_log_force[7301] <= 1'h0;
      write_enable_data_log_force[7302] <= 1'h0;
      write_enable_data_log_force[7303] <= 1'h0;
      write_enable_data_log_force[7304] <= 1'h0;
      write_enable_data_log_force[7305] <= 1'h0;
      write_enable_data_log_force[7306] <= 1'h0;
      write_enable_data_log_force[7307] <= 1'h0;
      write_enable_data_log_force[7308] <= 1'h0;
      write_enable_data_log_force[7309] <= 1'h0;
      write_enable_data_log_force[7310] <= 1'h0;
      write_enable_data_log_force[7311] <= 1'h0;
      write_enable_data_log_force[7312] <= 1'h0;
      write_enable_data_log_force[7313] <= 1'h0;
      write_enable_data_log_force[7314] <= 1'h0;
      write_enable_data_log_force[7315] <= 1'h0;
      write_enable_data_log_force[7316] <= 1'h0;
      write_enable_data_log_force[7317] <= 1'h0;
      write_enable_data_log_force[7318] <= 1'h0;
      write_enable_data_log_force[7319] <= 1'h0;
      write_enable_data_log_force[7320] <= 1'h0;
      write_enable_data_log_force[7321] <= 1'h0;
      write_enable_data_log_force[7322] <= 1'h0;
      write_enable_data_log_force[7323] <= 1'h0;
      write_enable_data_log_force[7324] <= 1'h0;
      write_enable_data_log_force[7325] <= 1'h0;
      write_enable_data_log_force[7326] <= 1'h0;
      write_enable_data_log_force[7327] <= 1'h0;
      write_enable_data_log_force[7328] <= 1'h0;
      write_enable_data_log_force[7329] <= 1'h0;
      write_enable_data_log_force[7330] <= 1'h0;
      write_enable_data_log_force[7331] <= 1'h0;
      write_enable_data_log_force[7332] <= 1'h0;
      write_enable_data_log_force[7333] <= 1'h0;
      write_enable_data_log_force[7334] <= 1'h0;
      write_enable_data_log_force[7335] <= 1'h0;
      write_enable_data_log_force[7336] <= 1'h0;
      write_enable_data_log_force[7337] <= 1'h0;
      write_enable_data_log_force[7338] <= 1'h0;
      write_enable_data_log_force[7339] <= 1'h0;
      write_enable_data_log_force[7340] <= 1'h0;
      write_enable_data_log_force[7341] <= 1'h0;
      write_enable_data_log_force[7342] <= 1'h0;
      write_enable_data_log_force[7343] <= 1'h0;
      write_enable_data_log_force[7344] <= 1'h0;
      write_enable_data_log_force[7345] <= 1'h0;
      write_enable_data_log_force[7346] <= 1'h0;
      write_enable_data_log_force[7347] <= 1'h0;
      write_enable_data_log_force[7348] <= 1'h0;
      write_enable_data_log_force[7349] <= 1'h0;
      write_enable_data_log_force[7350] <= 1'h0;
      write_enable_data_log_force[7351] <= 1'h0;
      write_enable_data_log_force[7352] <= 1'h0;
      write_enable_data_log_force[7353] <= 1'h0;
      write_enable_data_log_force[7354] <= 1'h0;
      write_enable_data_log_force[7355] <= 1'h0;
      write_enable_data_log_force[7356] <= 1'h0;
      write_enable_data_log_force[7357] <= 1'h0;
      write_enable_data_log_force[7358] <= 1'h0;
      write_enable_data_log_force[7359] <= 1'h0;
      write_enable_data_log_force[7360] <= 1'h0;
      write_enable_data_log_force[7361] <= 1'h0;
      write_enable_data_log_force[7362] <= 1'h0;
      write_enable_data_log_force[7363] <= 1'h0;
      write_enable_data_log_force[7364] <= 1'h0;
      write_enable_data_log_force[7365] <= 1'h0;
      write_enable_data_log_force[7366] <= 1'h0;
      write_enable_data_log_force[7367] <= 1'h0;
      write_enable_data_log_force[7368] <= 1'h0;
      write_enable_data_log_force[7369] <= 1'h0;
      write_enable_data_log_force[7370] <= 1'h0;
      write_enable_data_log_force[7371] <= 1'h0;
      write_enable_data_log_force[7372] <= 1'h0;
      write_enable_data_log_force[7373] <= 1'h0;
      write_enable_data_log_force[7374] <= 1'h0;
      write_enable_data_log_force[7375] <= 1'h0;
      write_enable_data_log_force[7376] <= 1'h0;
      write_enable_data_log_force[7377] <= 1'h0;
      write_enable_data_log_force[7378] <= 1'h0;
      write_enable_data_log_force[7379] <= 1'h0;
      write_enable_data_log_force[7380] <= 1'h0;
      write_enable_data_log_force[7381] <= 1'h0;
      write_enable_data_log_force[7382] <= 1'h0;
      write_enable_data_log_force[7383] <= 1'h0;
      write_enable_data_log_force[7384] <= 1'h0;
      write_enable_data_log_force[7385] <= 1'h0;
      write_enable_data_log_force[7386] <= 1'h0;
      write_enable_data_log_force[7387] <= 1'h0;
      write_enable_data_log_force[7388] <= 1'h0;
      write_enable_data_log_force[7389] <= 1'h0;
      write_enable_data_log_force[7390] <= 1'h0;
      write_enable_data_log_force[7391] <= 1'h0;
      write_enable_data_log_force[7392] <= 1'h0;
      write_enable_data_log_force[7393] <= 1'h0;
      write_enable_data_log_force[7394] <= 1'h0;
      write_enable_data_log_force[7395] <= 1'h0;
      write_enable_data_log_force[7396] <= 1'h0;
      write_enable_data_log_force[7397] <= 1'h0;
      write_enable_data_log_force[7398] <= 1'h0;
      write_enable_data_log_force[7399] <= 1'h0;
      write_enable_data_log_force[7400] <= 1'h0;
      write_enable_data_log_force[7401] <= 1'h0;
      write_enable_data_log_force[7402] <= 1'h0;
      write_enable_data_log_force[7403] <= 1'h0;
      write_enable_data_log_force[7404] <= 1'h0;
      write_enable_data_log_force[7405] <= 1'h0;
      write_enable_data_log_force[7406] <= 1'h0;
      write_enable_data_log_force[7407] <= 1'h0;
      write_enable_data_log_force[7408] <= 1'h0;
      write_enable_data_log_force[7409] <= 1'h0;
      write_enable_data_log_force[7410] <= 1'h0;
      write_enable_data_log_force[7411] <= 1'h0;
      write_enable_data_log_force[7412] <= 1'h0;
      write_enable_data_log_force[7413] <= 1'h0;
      write_enable_data_log_force[7414] <= 1'h0;
      write_enable_data_log_force[7415] <= 1'h0;
      write_enable_data_log_force[7416] <= 1'h0;
      write_enable_data_log_force[7417] <= 1'h0;
      write_enable_data_log_force[7418] <= 1'h0;
      write_enable_data_log_force[7419] <= 1'h0;
      write_enable_data_log_force[7420] <= 1'h0;
      write_enable_data_log_force[7421] <= 1'h0;
      write_enable_data_log_force[7422] <= 1'h0;
      write_enable_data_log_force[7423] <= 1'h0;
      write_enable_data_log_force[7424] <= 1'h0;
      write_enable_data_log_force[7425] <= 1'h0;
      write_enable_data_log_force[7426] <= 1'h0;
      write_enable_data_log_force[7427] <= 1'h0;
      write_enable_data_log_force[7428] <= 1'h0;
      write_enable_data_log_force[7429] <= 1'h0;
      write_enable_data_log_force[7430] <= 1'h0;
      write_enable_data_log_force[7431] <= 1'h0;
      write_enable_data_log_force[7432] <= 1'h0;
      write_enable_data_log_force[7433] <= 1'h0;
      write_enable_data_log_force[7434] <= 1'h0;
      write_enable_data_log_force[7435] <= 1'h0;
      write_enable_data_log_force[7436] <= 1'h0;
      write_enable_data_log_force[7437] <= 1'h0;
      write_enable_data_log_force[7438] <= 1'h0;
      write_enable_data_log_force[7439] <= 1'h0;
      write_enable_data_log_force[7440] <= 1'h0;
      write_enable_data_log_force[7441] <= 1'h0;
      write_enable_data_log_force[7442] <= 1'h0;
      write_enable_data_log_force[7443] <= 1'h0;
      write_enable_data_log_force[7444] <= 1'h0;
      write_enable_data_log_force[7445] <= 1'h0;
      write_enable_data_log_force[7446] <= 1'h0;
      write_enable_data_log_force[7447] <= 1'h0;
      write_enable_data_log_force[7448] <= 1'h0;
      write_enable_data_log_force[7449] <= 1'h0;
      write_enable_data_log_force[7450] <= 1'h0;
      write_enable_data_log_force[7451] <= 1'h0;
      write_enable_data_log_force[7452] <= 1'h0;
      write_enable_data_log_force[7453] <= 1'h0;
      write_enable_data_log_force[7454] <= 1'h0;
      write_enable_data_log_force[7455] <= 1'h0;
      write_enable_data_log_force[7456] <= 1'h0;
      write_enable_data_log_force[7457] <= 1'h0;
      write_enable_data_log_force[7458] <= 1'h0;
      write_enable_data_log_force[7459] <= 1'h0;
      write_enable_data_log_force[7460] <= 1'h0;
      write_enable_data_log_force[7461] <= 1'h0;
      write_enable_data_log_force[7462] <= 1'h0;
      write_enable_data_log_force[7463] <= 1'h0;
      write_enable_data_log_force[7464] <= 1'h0;
      write_enable_data_log_force[7465] <= 1'h0;
      write_enable_data_log_force[7466] <= 1'h0;
      write_enable_data_log_force[7467] <= 1'h0;
      write_enable_data_log_force[7468] <= 1'h0;
      write_enable_data_log_force[7469] <= 1'h0;
      write_enable_data_log_force[7470] <= 1'h0;
      write_enable_data_log_force[7471] <= 1'h0;
      write_enable_data_log_force[7472] <= 1'h0;
      write_enable_data_log_force[7473] <= 1'h0;
      write_enable_data_log_force[7474] <= 1'h0;
      write_enable_data_log_force[7475] <= 1'h0;
      write_enable_data_log_force[7476] <= 1'h0;
      write_enable_data_log_force[7477] <= 1'h0;
      write_enable_data_log_force[7478] <= 1'h0;
      write_enable_data_log_force[7479] <= 1'h0;
      write_enable_data_log_force[7480] <= 1'h0;
      write_enable_data_log_force[7481] <= 1'h0;
      write_enable_data_log_force[7482] <= 1'h0;
      write_enable_data_log_force[7483] <= 1'h0;
      write_enable_data_log_force[7484] <= 1'h0;
      write_enable_data_log_force[7485] <= 1'h0;
      write_enable_data_log_force[7486] <= 1'h0;
      write_enable_data_log_force[7487] <= 1'h0;
      write_enable_data_log_force[7488] <= 1'h0;
      write_enable_data_log_force[7489] <= 1'h0;
      write_enable_data_log_force[7490] <= 1'h0;
      write_enable_data_log_force[7491] <= 1'h0;
      write_enable_data_log_force[7492] <= 1'h0;
      write_enable_data_log_force[7493] <= 1'h0;
      write_enable_data_log_force[7494] <= 1'h0;
      write_enable_data_log_force[7495] <= 1'h0;
      write_enable_data_log_force[7496] <= 1'h0;
      write_enable_data_log_force[7497] <= 1'h0;
      write_enable_data_log_force[7498] <= 1'h0;
      write_enable_data_log_force[7499] <= 1'h0;
      write_enable_data_log_force[7500] <= 1'h0;
      write_enable_data_log_force[7501] <= 1'h0;
      write_enable_data_log_force[7502] <= 1'h0;
      write_enable_data_log_force[7503] <= 1'h0;
      write_enable_data_log_force[7504] <= 1'h0;
      write_enable_data_log_force[7505] <= 1'h0;
      write_enable_data_log_force[7506] <= 1'h0;
      write_enable_data_log_force[7507] <= 1'h0;
      write_enable_data_log_force[7508] <= 1'h0;
      write_enable_data_log_force[7509] <= 1'h0;
      write_enable_data_log_force[7510] <= 1'h0;
      write_enable_data_log_force[7511] <= 1'h0;
      write_enable_data_log_force[7512] <= 1'h0;
      write_enable_data_log_force[7513] <= 1'h0;
      write_enable_data_log_force[7514] <= 1'h0;
      write_enable_data_log_force[7515] <= 1'h0;
      write_enable_data_log_force[7516] <= 1'h0;
      write_enable_data_log_force[7517] <= 1'h0;
      write_enable_data_log_force[7518] <= 1'h0;
      write_enable_data_log_force[7519] <= 1'h0;
      write_enable_data_log_force[7520] <= 1'h0;
      write_enable_data_log_force[7521] <= 1'h0;
      write_enable_data_log_force[7522] <= 1'h0;
      write_enable_data_log_force[7523] <= 1'h0;
      write_enable_data_log_force[7524] <= 1'h0;
      write_enable_data_log_force[7525] <= 1'h0;
      write_enable_data_log_force[7526] <= 1'h0;
      write_enable_data_log_force[7527] <= 1'h0;
      write_enable_data_log_force[7528] <= 1'h0;
      write_enable_data_log_force[7529] <= 1'h0;
      write_enable_data_log_force[7530] <= 1'h0;
      write_enable_data_log_force[7531] <= 1'h0;
      write_enable_data_log_force[7532] <= 1'h0;
      write_enable_data_log_force[7533] <= 1'h0;
      write_enable_data_log_force[7534] <= 1'h0;
      write_enable_data_log_force[7535] <= 1'h0;
      write_enable_data_log_force[7536] <= 1'h0;
      write_enable_data_log_force[7537] <= 1'h0;
      write_enable_data_log_force[7538] <= 1'h0;
      write_enable_data_log_force[7539] <= 1'h0;
      write_enable_data_log_force[7540] <= 1'h0;
      write_enable_data_log_force[7541] <= 1'h0;
      write_enable_data_log_force[7542] <= 1'h0;
      write_enable_data_log_force[7543] <= 1'h0;
      write_enable_data_log_force[7544] <= 1'h0;
      write_enable_data_log_force[7545] <= 1'h0;
      write_enable_data_log_force[7546] <= 1'h0;
      write_enable_data_log_force[7547] <= 1'h0;
      write_enable_data_log_force[7548] <= 1'h0;
      write_enable_data_log_force[7549] <= 1'h0;
      write_enable_data_log_force[7550] <= 1'h0;
      write_enable_data_log_force[7551] <= 1'h0;
      write_enable_data_log_force[7552] <= 1'h0;
      write_enable_data_log_force[7553] <= 1'h0;
      write_enable_data_log_force[7554] <= 1'h0;
      write_enable_data_log_force[7555] <= 1'h0;
      write_enable_data_log_force[7556] <= 1'h0;
      write_enable_data_log_force[7557] <= 1'h0;
      write_enable_data_log_force[7558] <= 1'h0;
      write_enable_data_log_force[7559] <= 1'h0;
      write_enable_data_log_force[7560] <= 1'h0;
      write_enable_data_log_force[7561] <= 1'h0;
      write_enable_data_log_force[7562] <= 1'h0;
      write_enable_data_log_force[7563] <= 1'h0;
      write_enable_data_log_force[7564] <= 1'h0;
      write_enable_data_log_force[7565] <= 1'h0;
      write_enable_data_log_force[7566] <= 1'h0;
      write_enable_data_log_force[7567] <= 1'h0;
      write_enable_data_log_force[7568] <= 1'h0;
      write_enable_data_log_force[7569] <= 1'h0;
      write_enable_data_log_force[7570] <= 1'h0;
      write_enable_data_log_force[7571] <= 1'h0;
      write_enable_data_log_force[7572] <= 1'h0;
      write_enable_data_log_force[7573] <= 1'h0;
      write_enable_data_log_force[7574] <= 1'h0;
      write_enable_data_log_force[7575] <= 1'h0;
      write_enable_data_log_force[7576] <= 1'h0;
      write_enable_data_log_force[7577] <= 1'h0;
      write_enable_data_log_force[7578] <= 1'h0;
      write_enable_data_log_force[7579] <= 1'h0;
      write_enable_data_log_force[7580] <= 1'h0;
      write_enable_data_log_force[7581] <= 1'h0;
      write_enable_data_log_force[7582] <= 1'h0;
      write_enable_data_log_force[7583] <= 1'h0;
      write_enable_data_log_force[7584] <= 1'h0;
      write_enable_data_log_force[7585] <= 1'h0;
      write_enable_data_log_force[7586] <= 1'h0;
      write_enable_data_log_force[7587] <= 1'h0;
      write_enable_data_log_force[7588] <= 1'h0;
      write_enable_data_log_force[7589] <= 1'h0;
      write_enable_data_log_force[7590] <= 1'h0;
      write_enable_data_log_force[7591] <= 1'h0;
      write_enable_data_log_force[7592] <= 1'h0;
      write_enable_data_log_force[7593] <= 1'h0;
      write_enable_data_log_force[7594] <= 1'h0;
      write_enable_data_log_force[7595] <= 1'h0;
      write_enable_data_log_force[7596] <= 1'h0;
      write_enable_data_log_force[7597] <= 1'h0;
      write_enable_data_log_force[7598] <= 1'h0;
      write_enable_data_log_force[7599] <= 1'h0;
      write_enable_data_log_force[7600] <= 1'h0;
      write_enable_data_log_force[7601] <= 1'h0;
      write_enable_data_log_force[7602] <= 1'h0;
      write_enable_data_log_force[7603] <= 1'h0;
      write_enable_data_log_force[7604] <= 1'h0;
      write_enable_data_log_force[7605] <= 1'h0;
      write_enable_data_log_force[7606] <= 1'h0;
      write_enable_data_log_force[7607] <= 1'h0;
      write_enable_data_log_force[7608] <= 1'h0;
      write_enable_data_log_force[7609] <= 1'h0;
      write_enable_data_log_force[7610] <= 1'h0;
      write_enable_data_log_force[7611] <= 1'h0;
      write_enable_data_log_force[7612] <= 1'h0;
      write_enable_data_log_force[7613] <= 1'h0;
      write_enable_data_log_force[7614] <= 1'h0;
      write_enable_data_log_force[7615] <= 1'h0;
      write_enable_data_log_force[7616] <= 1'h0;
      write_enable_data_log_force[7617] <= 1'h0;
      write_enable_data_log_force[7618] <= 1'h0;
      write_enable_data_log_force[7619] <= 1'h0;
      write_enable_data_log_force[7620] <= 1'h0;
      write_enable_data_log_force[7621] <= 1'h0;
      write_enable_data_log_force[7622] <= 1'h0;
      write_enable_data_log_force[7623] <= 1'h0;
      write_enable_data_log_force[7624] <= 1'h0;
      write_enable_data_log_force[7625] <= 1'h0;
      write_enable_data_log_force[7626] <= 1'h0;
      write_enable_data_log_force[7627] <= 1'h0;
      write_enable_data_log_force[7628] <= 1'h0;
      write_enable_data_log_force[7629] <= 1'h0;
      write_enable_data_log_force[7630] <= 1'h0;
      write_enable_data_log_force[7631] <= 1'h0;
      write_enable_data_log_force[7632] <= 1'h0;
      write_enable_data_log_force[7633] <= 1'h0;
      write_enable_data_log_force[7634] <= 1'h0;
      write_enable_data_log_force[7635] <= 1'h0;
      write_enable_data_log_force[7636] <= 1'h0;
      write_enable_data_log_force[7637] <= 1'h0;
      write_enable_data_log_force[7638] <= 1'h0;
      write_enable_data_log_force[7639] <= 1'h0;
      write_enable_data_log_force[7640] <= 1'h0;
      write_enable_data_log_force[7641] <= 1'h0;
      write_enable_data_log_force[7642] <= 1'h0;
      write_enable_data_log_force[7643] <= 1'h0;
      write_enable_data_log_force[7644] <= 1'h0;
      write_enable_data_log_force[7645] <= 1'h0;
      write_enable_data_log_force[7646] <= 1'h0;
      write_enable_data_log_force[7647] <= 1'h0;
      write_enable_data_log_force[7648] <= 1'h0;
      write_enable_data_log_force[7649] <= 1'h0;
      write_enable_data_log_force[7650] <= 1'h0;
      write_enable_data_log_force[7651] <= 1'h0;
      write_enable_data_log_force[7652] <= 1'h0;
      write_enable_data_log_force[7653] <= 1'h0;
      write_enable_data_log_force[7654] <= 1'h0;
      write_enable_data_log_force[7655] <= 1'h0;
      write_enable_data_log_force[7656] <= 1'h0;
      write_enable_data_log_force[7657] <= 1'h0;
      write_enable_data_log_force[7658] <= 1'h0;
      write_enable_data_log_force[7659] <= 1'h0;
      write_enable_data_log_force[7660] <= 1'h0;
      write_enable_data_log_force[7661] <= 1'h0;
      write_enable_data_log_force[7662] <= 1'h0;
      write_enable_data_log_force[7663] <= 1'h0;
      write_enable_data_log_force[7664] <= 1'h0;
      write_enable_data_log_force[7665] <= 1'h0;
      write_enable_data_log_force[7666] <= 1'h0;
      write_enable_data_log_force[7667] <= 1'h0;
      write_enable_data_log_force[7668] <= 1'h0;
      write_enable_data_log_force[7669] <= 1'h0;
      write_enable_data_log_force[7670] <= 1'h0;
      write_enable_data_log_force[7671] <= 1'h0;
      write_enable_data_log_force[7672] <= 1'h0;
      write_enable_data_log_force[7673] <= 1'h0;
      write_enable_data_log_force[7674] <= 1'h0;
      write_enable_data_log_force[7675] <= 1'h0;
      write_enable_data_log_force[7676] <= 1'h0;
      write_enable_data_log_force[7677] <= 1'h0;
      write_enable_data_log_force[7678] <= 1'h0;
      write_enable_data_log_force[7679] <= 1'h0;
      write_enable_data_log_force[7680] <= 1'h0;
      write_enable_data_log_force[7681] <= 1'h0;
      write_enable_data_log_force[7682] <= 1'h0;
      write_enable_data_log_force[7683] <= 1'h0;
      write_enable_data_log_force[7684] <= 1'h0;
      write_enable_data_log_force[7685] <= 1'h0;
      write_enable_data_log_force[7686] <= 1'h0;
      write_enable_data_log_force[7687] <= 1'h0;
      write_enable_data_log_force[7688] <= 1'h0;
      write_enable_data_log_force[7689] <= 1'h0;
      write_enable_data_log_force[7690] <= 1'h0;
      write_enable_data_log_force[7691] <= 1'h0;
      write_enable_data_log_force[7692] <= 1'h0;
      write_enable_data_log_force[7693] <= 1'h0;
      write_enable_data_log_force[7694] <= 1'h0;
      write_enable_data_log_force[7695] <= 1'h0;
      write_enable_data_log_force[7696] <= 1'h0;
      write_enable_data_log_force[7697] <= 1'h0;
      write_enable_data_log_force[7698] <= 1'h0;
      write_enable_data_log_force[7699] <= 1'h0;
      write_enable_data_log_force[7700] <= 1'h0;
      write_enable_data_log_force[7701] <= 1'h0;
      write_enable_data_log_force[7702] <= 1'h0;
      write_enable_data_log_force[7703] <= 1'h0;
      write_enable_data_log_force[7704] <= 1'h0;
      write_enable_data_log_force[7705] <= 1'h0;
      write_enable_data_log_force[7706] <= 1'h0;
      write_enable_data_log_force[7707] <= 1'h0;
      write_enable_data_log_force[7708] <= 1'h0;
      write_enable_data_log_force[7709] <= 1'h0;
      write_enable_data_log_force[7710] <= 1'h0;
      write_enable_data_log_force[7711] <= 1'h0;
      write_enable_data_log_force[7712] <= 1'h0;
      write_enable_data_log_force[7713] <= 1'h0;
      write_enable_data_log_force[7714] <= 1'h0;
      write_enable_data_log_force[7715] <= 1'h0;
      write_enable_data_log_force[7716] <= 1'h0;
      write_enable_data_log_force[7717] <= 1'h0;
      write_enable_data_log_force[7718] <= 1'h0;
      write_enable_data_log_force[7719] <= 1'h0;
      write_enable_data_log_force[7720] <= 1'h0;
      write_enable_data_log_force[7721] <= 1'h0;
      write_enable_data_log_force[7722] <= 1'h0;
      write_enable_data_log_force[7723] <= 1'h0;
      write_enable_data_log_force[7724] <= 1'h0;
      write_enable_data_log_force[7725] <= 1'h0;
      write_enable_data_log_force[7726] <= 1'h0;
      write_enable_data_log_force[7727] <= 1'h0;
      write_enable_data_log_force[7728] <= 1'h0;
      write_enable_data_log_force[7729] <= 1'h0;
      write_enable_data_log_force[7730] <= 1'h0;
      write_enable_data_log_force[7731] <= 1'h0;
      write_enable_data_log_force[7732] <= 1'h0;
      write_enable_data_log_force[7733] <= 1'h0;
      write_enable_data_log_force[7734] <= 1'h0;
      write_enable_data_log_force[7735] <= 1'h0;
      write_enable_data_log_force[7736] <= 1'h0;
      write_enable_data_log_force[7737] <= 1'h0;
      write_enable_data_log_force[7738] <= 1'h0;
      write_enable_data_log_force[7739] <= 1'h0;
      write_enable_data_log_force[7740] <= 1'h0;
      write_enable_data_log_force[7741] <= 1'h0;
      write_enable_data_log_force[7742] <= 1'h0;
      write_enable_data_log_force[7743] <= 1'h0;
      write_enable_data_log_force[7744] <= 1'h0;
      write_enable_data_log_force[7745] <= 1'h0;
      write_enable_data_log_force[7746] <= 1'h0;
      write_enable_data_log_force[7747] <= 1'h0;
      write_enable_data_log_force[7748] <= 1'h0;
      write_enable_data_log_force[7749] <= 1'h0;
      write_enable_data_log_force[7750] <= 1'h0;
      write_enable_data_log_force[7751] <= 1'h0;
      write_enable_data_log_force[7752] <= 1'h0;
      write_enable_data_log_force[7753] <= 1'h0;
      write_enable_data_log_force[7754] <= 1'h0;
      write_enable_data_log_force[7755] <= 1'h0;
      write_enable_data_log_force[7756] <= 1'h0;
      write_enable_data_log_force[7757] <= 1'h0;
      write_enable_data_log_force[7758] <= 1'h0;
      write_enable_data_log_force[7759] <= 1'h0;
      write_enable_data_log_force[7760] <= 1'h0;
      write_enable_data_log_force[7761] <= 1'h0;
      write_enable_data_log_force[7762] <= 1'h0;
      write_enable_data_log_force[7763] <= 1'h0;
      write_enable_data_log_force[7764] <= 1'h0;
      write_enable_data_log_force[7765] <= 1'h0;
      write_enable_data_log_force[7766] <= 1'h0;
      write_enable_data_log_force[7767] <= 1'h0;
      write_enable_data_log_force[7768] <= 1'h0;
      write_enable_data_log_force[7769] <= 1'h0;
      write_enable_data_log_force[7770] <= 1'h0;
      write_enable_data_log_force[7771] <= 1'h0;
      write_enable_data_log_force[7772] <= 1'h0;
      write_enable_data_log_force[7773] <= 1'h0;
      write_enable_data_log_force[7774] <= 1'h0;
      write_enable_data_log_force[7775] <= 1'h0;
      write_enable_data_log_force[7776] <= 1'h0;
      write_enable_data_log_force[7777] <= 1'h0;
      write_enable_data_log_force[7778] <= 1'h0;
      write_enable_data_log_force[7779] <= 1'h0;
      write_enable_data_log_force[7780] <= 1'h0;
      write_enable_data_log_force[7781] <= 1'h0;
      write_enable_data_log_force[7782] <= 1'h0;
      write_enable_data_log_force[7783] <= 1'h0;
      write_enable_data_log_force[7784] <= 1'h0;
      write_enable_data_log_force[7785] <= 1'h0;
      write_enable_data_log_force[7786] <= 1'h0;
      write_enable_data_log_force[7787] <= 1'h0;
      write_enable_data_log_force[7788] <= 1'h0;
      write_enable_data_log_force[7789] <= 1'h0;
      write_enable_data_log_force[7790] <= 1'h0;
      write_enable_data_log_force[7791] <= 1'h0;
      write_enable_data_log_force[7792] <= 1'h0;
      write_enable_data_log_force[7793] <= 1'h0;
      write_enable_data_log_force[7794] <= 1'h0;
      write_enable_data_log_force[7795] <= 1'h0;
      write_enable_data_log_force[7796] <= 1'h0;
      write_enable_data_log_force[7797] <= 1'h0;
      write_enable_data_log_force[7798] <= 1'h0;
      write_enable_data_log_force[7799] <= 1'h0;
      write_enable_data_log_force[7800] <= 1'h0;
      write_enable_data_log_force[7801] <= 1'h0;
      write_enable_data_log_force[7802] <= 1'h0;
      write_enable_data_log_force[7803] <= 1'h0;
      write_enable_data_log_force[7804] <= 1'h0;
      write_enable_data_log_force[7805] <= 1'h0;
      write_enable_data_log_force[7806] <= 1'h0;
      write_enable_data_log_force[7807] <= 1'h0;
      write_enable_data_log_force[7808] <= 1'h0;
      write_enable_data_log_force[7809] <= 1'h0;
      write_enable_data_log_force[7810] <= 1'h0;
      write_enable_data_log_force[7811] <= 1'h0;
      write_enable_data_log_force[7812] <= 1'h0;
      write_enable_data_log_force[7813] <= 1'h0;
      write_enable_data_log_force[7814] <= 1'h0;
      write_enable_data_log_force[7815] <= 1'h0;
      write_enable_data_log_force[7816] <= 1'h0;
      write_enable_data_log_force[7817] <= 1'h0;
      write_enable_data_log_force[7818] <= 1'h0;
      write_enable_data_log_force[7819] <= 1'h0;
      write_enable_data_log_force[7820] <= 1'h0;
      write_enable_data_log_force[7821] <= 1'h0;
      write_enable_data_log_force[7822] <= 1'h0;
      write_enable_data_log_force[7823] <= 1'h0;
      write_enable_data_log_force[7824] <= 1'h0;
      write_enable_data_log_force[7825] <= 1'h0;
      write_enable_data_log_force[7826] <= 1'h0;
      write_enable_data_log_force[7827] <= 1'h0;
      write_enable_data_log_force[7828] <= 1'h0;
      write_enable_data_log_force[7829] <= 1'h0;
      write_enable_data_log_force[7830] <= 1'h0;
      write_enable_data_log_force[7831] <= 1'h0;
      write_enable_data_log_force[7832] <= 1'h0;
      write_enable_data_log_force[7833] <= 1'h0;
      write_enable_data_log_force[7834] <= 1'h0;
      write_enable_data_log_force[7835] <= 1'h0;
      write_enable_data_log_force[7836] <= 1'h0;
      write_enable_data_log_force[7837] <= 1'h0;
      write_enable_data_log_force[7838] <= 1'h0;
      write_enable_data_log_force[7839] <= 1'h0;
      write_enable_data_log_force[7840] <= 1'h0;
      write_enable_data_log_force[7841] <= 1'h0;
      write_enable_data_log_force[7842] <= 1'h0;
      write_enable_data_log_force[7843] <= 1'h0;
      write_enable_data_log_force[7844] <= 1'h0;
      write_enable_data_log_force[7845] <= 1'h0;
      write_enable_data_log_force[7846] <= 1'h0;
      write_enable_data_log_force[7847] <= 1'h0;
      write_enable_data_log_force[7848] <= 1'h0;
      write_enable_data_log_force[7849] <= 1'h0;
      write_enable_data_log_force[7850] <= 1'h0;
      write_enable_data_log_force[7851] <= 1'h0;
      write_enable_data_log_force[7852] <= 1'h0;
      write_enable_data_log_force[7853] <= 1'h0;
      write_enable_data_log_force[7854] <= 1'h0;
      write_enable_data_log_force[7855] <= 1'h0;
      write_enable_data_log_force[7856] <= 1'h0;
      write_enable_data_log_force[7857] <= 1'h0;
      write_enable_data_log_force[7858] <= 1'h0;
      write_enable_data_log_force[7859] <= 1'h0;
      write_enable_data_log_force[7860] <= 1'h0;
      write_enable_data_log_force[7861] <= 1'h0;
      write_enable_data_log_force[7862] <= 1'h0;
      write_enable_data_log_force[7863] <= 1'h0;
      write_enable_data_log_force[7864] <= 1'h0;
      write_enable_data_log_force[7865] <= 1'h0;
      write_enable_data_log_force[7866] <= 1'h0;
      write_enable_data_log_force[7867] <= 1'h0;
      write_enable_data_log_force[7868] <= 1'h0;
      write_enable_data_log_force[7869] <= 1'h0;
      write_enable_data_log_force[7870] <= 1'h0;
      write_enable_data_log_force[7871] <= 1'h0;
      write_enable_data_log_force[7872] <= 1'h0;
      write_enable_data_log_force[7873] <= 1'h0;
      write_enable_data_log_force[7874] <= 1'h0;
      write_enable_data_log_force[7875] <= 1'h0;
      write_enable_data_log_force[7876] <= 1'h0;
      write_enable_data_log_force[7877] <= 1'h0;
      write_enable_data_log_force[7878] <= 1'h0;
      write_enable_data_log_force[7879] <= 1'h0;
      write_enable_data_log_force[7880] <= 1'h0;
      write_enable_data_log_force[7881] <= 1'h0;
      write_enable_data_log_force[7882] <= 1'h0;
      write_enable_data_log_force[7883] <= 1'h0;
      write_enable_data_log_force[7884] <= 1'h0;
      write_enable_data_log_force[7885] <= 1'h0;
      write_enable_data_log_force[7886] <= 1'h0;
      write_enable_data_log_force[7887] <= 1'h0;
      write_enable_data_log_force[7888] <= 1'h0;
      write_enable_data_log_force[7889] <= 1'h0;
      write_enable_data_log_force[7890] <= 1'h0;
      write_enable_data_log_force[7891] <= 1'h0;
      write_enable_data_log_force[7892] <= 1'h0;
      write_enable_data_log_force[7893] <= 1'h0;
      write_enable_data_log_force[7894] <= 1'h0;
      write_enable_data_log_force[7895] <= 1'h0;
      write_enable_data_log_force[7896] <= 1'h0;
      write_enable_data_log_force[7897] <= 1'h0;
      write_enable_data_log_force[7898] <= 1'h0;
      write_enable_data_log_force[7899] <= 1'h0;
      write_enable_data_log_force[7900] <= 1'h0;
      write_enable_data_log_force[7901] <= 1'h0;
      write_enable_data_log_force[7902] <= 1'h0;
      write_enable_data_log_force[7903] <= 1'h0;
      write_enable_data_log_force[7904] <= 1'h0;
      write_enable_data_log_force[7905] <= 1'h0;
      write_enable_data_log_force[7906] <= 1'h0;
      write_enable_data_log_force[7907] <= 1'h0;
      write_enable_data_log_force[7908] <= 1'h0;
      write_enable_data_log_force[7909] <= 1'h0;
      write_enable_data_log_force[7910] <= 1'h0;
      write_enable_data_log_force[7911] <= 1'h0;
      write_enable_data_log_force[7912] <= 1'h0;
      write_enable_data_log_force[7913] <= 1'h0;
      write_enable_data_log_force[7914] <= 1'h0;
      write_enable_data_log_force[7915] <= 1'h0;
      write_enable_data_log_force[7916] <= 1'h0;
      write_enable_data_log_force[7917] <= 1'h0;
      write_enable_data_log_force[7918] <= 1'h0;
      write_enable_data_log_force[7919] <= 1'h0;
      write_enable_data_log_force[7920] <= 1'h0;
      write_enable_data_log_force[7921] <= 1'h0;
      write_enable_data_log_force[7922] <= 1'h0;
      write_enable_data_log_force[7923] <= 1'h0;
      write_enable_data_log_force[7924] <= 1'h0;
      write_enable_data_log_force[7925] <= 1'h0;
      write_enable_data_log_force[7926] <= 1'h0;
      write_enable_data_log_force[7927] <= 1'h0;
      write_enable_data_log_force[7928] <= 1'h0;
      write_enable_data_log_force[7929] <= 1'h0;
      write_enable_data_log_force[7930] <= 1'h0;
      write_enable_data_log_force[7931] <= 1'h0;
      write_enable_data_log_force[7932] <= 1'h0;
      write_enable_data_log_force[7933] <= 1'h0;
      write_enable_data_log_force[7934] <= 1'h0;
      write_enable_data_log_force[7935] <= 1'h0;
      write_enable_data_log_force[7936] <= 1'h0;
      write_enable_data_log_force[7937] <= 1'h0;
      write_enable_data_log_force[7938] <= 1'h0;
      write_enable_data_log_force[7939] <= 1'h0;
      write_enable_data_log_force[7940] <= 1'h0;
      write_enable_data_log_force[7941] <= 1'h0;
      write_enable_data_log_force[7942] <= 1'h0;
      write_enable_data_log_force[7943] <= 1'h0;
      write_enable_data_log_force[7944] <= 1'h0;
      write_enable_data_log_force[7945] <= 1'h0;
      write_enable_data_log_force[7946] <= 1'h0;
      write_enable_data_log_force[7947] <= 1'h0;
      write_enable_data_log_force[7948] <= 1'h0;
      write_enable_data_log_force[7949] <= 1'h0;
      write_enable_data_log_force[7950] <= 1'h0;
      write_enable_data_log_force[7951] <= 1'h0;
      write_enable_data_log_force[7952] <= 1'h0;
      write_enable_data_log_force[7953] <= 1'h0;
      write_enable_data_log_force[7954] <= 1'h0;
      write_enable_data_log_force[7955] <= 1'h0;
      write_enable_data_log_force[7956] <= 1'h0;
      write_enable_data_log_force[7957] <= 1'h0;
      write_enable_data_log_force[7958] <= 1'h0;
      write_enable_data_log_force[7959] <= 1'h0;
      write_enable_data_log_force[7960] <= 1'h0;
      write_enable_data_log_force[7961] <= 1'h0;
      write_enable_data_log_force[7962] <= 1'h0;
      write_enable_data_log_force[7963] <= 1'h0;
      write_enable_data_log_force[7964] <= 1'h0;
      write_enable_data_log_force[7965] <= 1'h0;
      write_enable_data_log_force[7966] <= 1'h0;
      write_enable_data_log_force[7967] <= 1'h0;
      write_enable_data_log_force[7968] <= 1'h0;
      write_enable_data_log_force[7969] <= 1'h0;
      write_enable_data_log_force[7970] <= 1'h0;
      write_enable_data_log_force[7971] <= 1'h0;
      write_enable_data_log_force[7972] <= 1'h0;
      write_enable_data_log_force[7973] <= 1'h0;
      write_enable_data_log_force[7974] <= 1'h0;
      write_enable_data_log_force[7975] <= 1'h0;
      write_enable_data_log_force[7976] <= 1'h0;
      write_enable_data_log_force[7977] <= 1'h0;
      write_enable_data_log_force[7978] <= 1'h0;
      write_enable_data_log_force[7979] <= 1'h0;
      write_enable_data_log_force[7980] <= 1'h0;
      write_enable_data_log_force[7981] <= 1'h0;
      write_enable_data_log_force[7982] <= 1'h0;
      write_enable_data_log_force[7983] <= 1'h0;
      write_enable_data_log_force[7984] <= 1'h0;
      write_enable_data_log_force[7985] <= 1'h0;
      write_enable_data_log_force[7986] <= 1'h0;
      write_enable_data_log_force[7987] <= 1'h0;
      write_enable_data_log_force[7988] <= 1'h0;
      write_enable_data_log_force[7989] <= 1'h0;
      write_enable_data_log_force[7990] <= 1'h0;
      write_enable_data_log_force[7991] <= 1'h0;
      write_enable_data_log_force[7992] <= 1'h0;
      write_enable_data_log_force[7993] <= 1'h0;
      write_enable_data_log_force[7994] <= 1'h0;
      write_enable_data_log_force[7995] <= 1'h0;
      write_enable_data_log_force[7996] <= 1'h0;
      write_enable_data_log_force[7997] <= 1'h0;
      write_enable_data_log_force[7998] <= 1'h0;
      write_enable_data_log_force[7999] <= 1'h0;
      write_enable_data_log_force[8000] <= 1'h0;
      write_enable_data_log_force[8001] <= 1'h0;
      write_enable_data_log_force[8002] <= 1'h0;
      write_enable_data_log_force[8003] <= 1'h0;
      write_enable_data_log_force[8004] <= 1'h0;
      write_enable_data_log_force[8005] <= 1'h0;
      write_enable_data_log_force[8006] <= 1'h0;
      write_enable_data_log_force[8007] <= 1'h0;
      write_enable_data_log_force[8008] <= 1'h0;
      write_enable_data_log_force[8009] <= 1'h0;
      write_enable_data_log_force[8010] <= 1'h0;
      write_enable_data_log_force[8011] <= 1'h0;
      write_enable_data_log_force[8012] <= 1'h0;
      write_enable_data_log_force[8013] <= 1'h0;
      write_enable_data_log_force[8014] <= 1'h0;
      write_enable_data_log_force[8015] <= 1'h0;
      write_enable_data_log_force[8016] <= 1'h0;
      write_enable_data_log_force[8017] <= 1'h0;
      write_enable_data_log_force[8018] <= 1'h0;
      write_enable_data_log_force[8019] <= 1'h0;
      write_enable_data_log_force[8020] <= 1'h0;
      write_enable_data_log_force[8021] <= 1'h0;
      write_enable_data_log_force[8022] <= 1'h0;
      write_enable_data_log_force[8023] <= 1'h0;
      write_enable_data_log_force[8024] <= 1'h0;
      write_enable_data_log_force[8025] <= 1'h0;
      write_enable_data_log_force[8026] <= 1'h0;
      write_enable_data_log_force[8027] <= 1'h0;
      write_enable_data_log_force[8028] <= 1'h0;
      write_enable_data_log_force[8029] <= 1'h0;
      write_enable_data_log_force[8030] <= 1'h0;
      write_enable_data_log_force[8031] <= 1'h0;
      write_enable_data_log_force[8032] <= 1'h0;
      write_enable_data_log_force[8033] <= 1'h0;
      write_enable_data_log_force[8034] <= 1'h0;
      write_enable_data_log_force[8035] <= 1'h0;
      write_enable_data_log_force[8036] <= 1'h0;
      write_enable_data_log_force[8037] <= 1'h0;
      write_enable_data_log_force[8038] <= 1'h0;
      write_enable_data_log_force[8039] <= 1'h0;
      write_enable_data_log_force[8040] <= 1'h0;
      write_enable_data_log_force[8041] <= 1'h0;
      write_enable_data_log_force[8042] <= 1'h0;
      write_enable_data_log_force[8043] <= 1'h0;
      write_enable_data_log_force[8044] <= 1'h0;
      write_enable_data_log_force[8045] <= 1'h0;
      write_enable_data_log_force[8046] <= 1'h0;
      write_enable_data_log_force[8047] <= 1'h0;
      write_enable_data_log_force[8048] <= 1'h0;
      write_enable_data_log_force[8049] <= 1'h0;
      write_enable_data_log_force[8050] <= 1'h0;
      write_enable_data_log_force[8051] <= 1'h0;
      write_enable_data_log_force[8052] <= 1'h0;
      write_enable_data_log_force[8053] <= 1'h0;
      write_enable_data_log_force[8054] <= 1'h0;
      write_enable_data_log_force[8055] <= 1'h0;
      write_enable_data_log_force[8056] <= 1'h0;
      write_enable_data_log_force[8057] <= 1'h0;
      write_enable_data_log_force[8058] <= 1'h0;
      write_enable_data_log_force[8059] <= 1'h0;
      write_enable_data_log_force[8060] <= 1'h0;
      write_enable_data_log_force[8061] <= 1'h0;
      write_enable_data_log_force[8062] <= 1'h0;
      write_enable_data_log_force[8063] <= 1'h0;
      write_enable_data_log_force[8064] <= 1'h0;
      write_enable_data_log_force[8065] <= 1'h0;
      write_enable_data_log_force[8066] <= 1'h0;
      write_enable_data_log_force[8067] <= 1'h0;
      write_enable_data_log_force[8068] <= 1'h0;
      write_enable_data_log_force[8069] <= 1'h0;
      write_enable_data_log_force[8070] <= 1'h0;
      write_enable_data_log_force[8071] <= 1'h0;
      write_enable_data_log_force[8072] <= 1'h0;
      write_enable_data_log_force[8073] <= 1'h0;
      write_enable_data_log_force[8074] <= 1'h0;
      write_enable_data_log_force[8075] <= 1'h0;
      write_enable_data_log_force[8076] <= 1'h0;
      write_enable_data_log_force[8077] <= 1'h0;
      write_enable_data_log_force[8078] <= 1'h0;
      write_enable_data_log_force[8079] <= 1'h0;
      write_enable_data_log_force[8080] <= 1'h0;
      write_enable_data_log_force[8081] <= 1'h0;
      write_enable_data_log_force[8082] <= 1'h0;
      write_enable_data_log_force[8083] <= 1'h0;
      write_enable_data_log_force[8084] <= 1'h0;
      write_enable_data_log_force[8085] <= 1'h0;
      write_enable_data_log_force[8086] <= 1'h0;
      write_enable_data_log_force[8087] <= 1'h0;
      write_enable_data_log_force[8088] <= 1'h0;
      write_enable_data_log_force[8089] <= 1'h0;
      write_enable_data_log_force[8090] <= 1'h0;
      write_enable_data_log_force[8091] <= 1'h0;
      write_enable_data_log_force[8092] <= 1'h0;
      write_enable_data_log_force[8093] <= 1'h0;
      write_enable_data_log_force[8094] <= 1'h0;
      write_enable_data_log_force[8095] <= 1'h0;
      write_enable_data_log_force[8096] <= 1'h0;
      write_enable_data_log_force[8097] <= 1'h0;
      write_enable_data_log_force[8098] <= 1'h0;
      write_enable_data_log_force[8099] <= 1'h0;
      write_enable_data_log_force[8100] <= 1'h0;
      write_enable_data_log_force[8101] <= 1'h0;
      write_enable_data_log_force[8102] <= 1'h0;
      write_enable_data_log_force[8103] <= 1'h0;
      write_enable_data_log_force[8104] <= 1'h0;
      write_enable_data_log_force[8105] <= 1'h0;
      write_enable_data_log_force[8106] <= 1'h0;
      write_enable_data_log_force[8107] <= 1'h0;
      write_enable_data_log_force[8108] <= 1'h0;
      write_enable_data_log_force[8109] <= 1'h0;
      write_enable_data_log_force[8110] <= 1'h0;
      write_enable_data_log_force[8111] <= 1'h0;
      write_enable_data_log_force[8112] <= 1'h0;
      write_enable_data_log_force[8113] <= 1'h0;
      write_enable_data_log_force[8114] <= 1'h0;
      write_enable_data_log_force[8115] <= 1'h0;
      write_enable_data_log_force[8116] <= 1'h0;
      write_enable_data_log_force[8117] <= 1'h0;
      write_enable_data_log_force[8118] <= 1'h0;
      write_enable_data_log_force[8119] <= 1'h0;
      write_enable_data_log_force[8120] <= 1'h0;
      write_enable_data_log_force[8121] <= 1'h0;
      write_enable_data_log_force[8122] <= 1'h0;
      write_enable_data_log_force[8123] <= 1'h0;
      write_enable_data_log_force[8124] <= 1'h0;
      write_enable_data_log_force[8125] <= 1'h0;
      write_enable_data_log_force[8126] <= 1'h0;
      write_enable_data_log_force[8127] <= 1'h0;
      write_enable_data_log_force[8128] <= 1'h0;
      write_enable_data_log_force[8129] <= 1'h0;
      write_enable_data_log_force[8130] <= 1'h0;
      write_enable_data_log_force[8131] <= 1'h0;
      write_enable_data_log_force[8132] <= 1'h0;
      write_enable_data_log_force[8133] <= 1'h0;
      write_enable_data_log_force[8134] <= 1'h0;
      write_enable_data_log_force[8135] <= 1'h0;
      write_enable_data_log_force[8136] <= 1'h0;
      write_enable_data_log_force[8137] <= 1'h0;
      write_enable_data_log_force[8138] <= 1'h0;
      write_enable_data_log_force[8139] <= 1'h0;
      write_enable_data_log_force[8140] <= 1'h0;
      write_enable_data_log_force[8141] <= 1'h0;
      write_enable_data_log_force[8142] <= 1'h0;
      write_enable_data_log_force[8143] <= 1'h0;
      write_enable_data_log_force[8144] <= 1'h0;
      write_enable_data_log_force[8145] <= 1'h0;
      write_enable_data_log_force[8146] <= 1'h0;
      write_enable_data_log_force[8147] <= 1'h0;
      write_enable_data_log_force[8148] <= 1'h0;
      write_enable_data_log_force[8149] <= 1'h0;
      write_enable_data_log_force[8150] <= 1'h0;
      write_enable_data_log_force[8151] <= 1'h0;
      write_enable_data_log_force[8152] <= 1'h0;
      write_enable_data_log_force[8153] <= 1'h0;
      write_enable_data_log_force[8154] <= 1'h0;
      write_enable_data_log_force[8155] <= 1'h0;
      write_enable_data_log_force[8156] <= 1'h0;
      write_enable_data_log_force[8157] <= 1'h0;
      write_enable_data_log_force[8158] <= 1'h0;
      write_enable_data_log_force[8159] <= 1'h0;
      write_enable_data_log_force[8160] <= 1'h0;
      write_enable_data_log_force[8161] <= 1'h0;
      write_enable_data_log_force[8162] <= 1'h0;
      write_enable_data_log_force[8163] <= 1'h0;
      write_enable_data_log_force[8164] <= 1'h0;
      write_enable_data_log_force[8165] <= 1'h0;
      write_enable_data_log_force[8166] <= 1'h0;
      write_enable_data_log_force[8167] <= 1'h0;
      write_enable_data_log_force[8168] <= 1'h0;
      write_enable_data_log_force[8169] <= 1'h0;
      write_enable_data_log_force[8170] <= 1'h0;
      write_enable_data_log_force[8171] <= 1'h0;
      write_enable_data_log_force[8172] <= 1'h0;
      write_enable_data_log_force[8173] <= 1'h0;
      write_enable_data_log_force[8174] <= 1'h0;
      write_enable_data_log_force[8175] <= 1'h0;
      write_enable_data_log_force[8176] <= 1'h0;
      write_enable_data_log_force[8177] <= 1'h0;
      write_enable_data_log_force[8178] <= 1'h0;
      write_enable_data_log_force[8179] <= 1'h0;
      write_enable_data_log_force[8180] <= 1'h0;
      write_enable_data_log_force[8181] <= 1'h0;
      write_enable_data_log_force[8182] <= 1'h0;
      write_enable_data_log_force[8183] <= 1'h0;
      write_enable_data_log_force[8184] <= 1'h0;
      write_enable_data_log_force[8185] <= 1'h0;
      write_enable_data_log_force[8186] <= 1'h0;
      write_enable_data_log_force[8187] <= 1'h0;
      write_enable_data_log_force[8188] <= 1'h0;
      write_enable_data_log_force[8189] <= 1'h0;
      write_enable_data_log_force[8190] <= 1'h0;
      write_enable_data_log_force[8191] <= 1'h0;
      write_enable_data_log_force[8192] <= 1'h0;
      write_enable_data_log_force[8193] <= 1'h0;
      write_enable_data_log_force[8194] <= 1'h0;
      write_enable_data_log_force[8195] <= 1'h0;
      write_enable_data_log_force[8196] <= 1'h0;
      write_enable_data_log_force[8197] <= 1'h0;
      write_enable_data_log_force[8198] <= 1'h0;
      write_enable_data_log_force[8199] <= 1'h0;
      write_enable_data_log_force[8200] <= 1'h0;
      write_enable_data_log_force[8201] <= 1'h0;
      write_enable_data_log_force[8202] <= 1'h0;
      write_enable_data_log_force[8203] <= 1'h0;
      write_enable_data_log_force[8204] <= 1'h0;
      write_enable_data_log_force[8205] <= 1'h0;
      write_enable_data_log_force[8206] <= 1'h0;
      write_enable_data_log_force[8207] <= 1'h0;
      write_enable_data_log_force[8208] <= 1'h0;
      write_enable_data_log_force[8209] <= 1'h0;
      write_enable_data_log_force[8210] <= 1'h0;
      write_enable_data_log_force[8211] <= 1'h0;
      write_enable_data_log_force[8212] <= 1'h0;
      write_enable_data_log_force[8213] <= 1'h0;
      write_enable_data_log_force[8214] <= 1'h0;
      write_enable_data_log_force[8215] <= 1'h0;
      write_enable_data_log_force[8216] <= 1'h0;
      write_enable_data_log_force[8217] <= 1'h0;
      write_enable_data_log_force[8218] <= 1'h0;
      write_enable_data_log_force[8219] <= 1'h0;
      write_enable_data_log_force[8220] <= 1'h0;
      write_enable_data_log_force[8221] <= 1'h0;
      write_enable_data_log_force[8222] <= 1'h0;
      write_enable_data_log_force[8223] <= 1'h0;
      write_enable_data_log_force[8224] <= 1'h0;
      write_enable_data_log_force[8225] <= 1'h0;
      write_enable_data_log_force[8226] <= 1'h0;
      write_enable_data_log_force[8227] <= 1'h0;
      write_enable_data_log_force[8228] <= 1'h0;
      write_enable_data_log_force[8229] <= 1'h0;
      write_enable_data_log_force[8230] <= 1'h0;
      write_enable_data_log_force[8231] <= 1'h0;
      write_enable_data_log_force[8232] <= 1'h0;
      write_enable_data_log_force[8233] <= 1'h0;
      write_enable_data_log_force[8234] <= 1'h0;
      write_enable_data_log_force[8235] <= 1'h0;
      write_enable_data_log_force[8236] <= 1'h0;
      write_enable_data_log_force[8237] <= 1'h0;
      write_enable_data_log_force[8238] <= 1'h0;
      write_enable_data_log_force[8239] <= 1'h0;
      write_enable_data_log_force[8240] <= 1'h0;
      write_enable_data_log_force[8241] <= 1'h0;
      write_enable_data_log_force[8242] <= 1'h0;
      write_enable_data_log_force[8243] <= 1'h0;
      write_enable_data_log_force[8244] <= 1'h0;
      write_enable_data_log_force[8245] <= 1'h0;
      write_enable_data_log_force[8246] <= 1'h0;
      write_enable_data_log_force[8247] <= 1'h0;
      write_enable_data_log_force[8248] <= 1'h0;
      write_enable_data_log_force[8249] <= 1'h0;
      write_enable_data_log_force[8250] <= 1'h0;
      write_enable_data_log_force[8251] <= 1'h0;
      write_enable_data_log_force[8252] <= 1'h0;
      write_enable_data_log_force[8253] <= 1'h0;
      write_enable_data_log_force[8254] <= 1'h0;
      write_enable_data_log_force[8255] <= 1'h0;
      write_enable_data_log_force[8256] <= 1'h0;
      write_enable_data_log_force[8257] <= 1'h0;
      write_enable_data_log_force[8258] <= 1'h0;
      write_enable_data_log_force[8259] <= 1'h0;
      write_enable_data_log_force[8260] <= 1'h0;
      write_enable_data_log_force[8261] <= 1'h0;
      write_enable_data_log_force[8262] <= 1'h0;
      write_enable_data_log_force[8263] <= 1'h0;
      write_enable_data_log_force[8264] <= 1'h0;
      write_enable_data_log_force[8265] <= 1'h0;
      write_enable_data_log_force[8266] <= 1'h0;
      write_enable_data_log_force[8267] <= 1'h0;
      write_enable_data_log_force[8268] <= 1'h0;
      write_enable_data_log_force[8269] <= 1'h0;
      write_enable_data_log_force[8270] <= 1'h0;
      write_enable_data_log_force[8271] <= 1'h0;
      write_enable_data_log_force[8272] <= 1'h0;
      write_enable_data_log_force[8273] <= 1'h0;
      write_enable_data_log_force[8274] <= 1'h0;
      write_enable_data_log_force[8275] <= 1'h0;
      write_enable_data_log_force[8276] <= 1'h0;
      write_enable_data_log_force[8277] <= 1'h0;
      write_enable_data_log_force[8278] <= 1'h0;
      write_enable_data_log_force[8279] <= 1'h0;
      write_enable_data_log_force[8280] <= 1'h0;
      write_enable_data_log_force[8281] <= 1'h0;
      write_enable_data_log_force[8282] <= 1'h0;
      write_enable_data_log_force[8283] <= 1'h0;
      write_enable_data_log_force[8284] <= 1'h0;
      write_enable_data_log_force[8285] <= 1'h0;
      write_enable_data_log_force[8286] <= 1'h0;
      write_enable_data_log_force[8287] <= 1'h0;
      write_enable_data_log_force[8288] <= 1'h0;
      write_enable_data_log_force[8289] <= 1'h0;
      write_enable_data_log_force[8290] <= 1'h0;
      write_enable_data_log_force[8291] <= 1'h0;
      write_enable_data_log_force[8292] <= 1'h0;
      write_enable_data_log_force[8293] <= 1'h0;
      write_enable_data_log_force[8294] <= 1'h0;
      write_enable_data_log_force[8295] <= 1'h0;
      write_enable_data_log_force[8296] <= 1'h0;
      write_enable_data_log_force[8297] <= 1'h0;
      write_enable_data_log_force[8298] <= 1'h0;
      write_enable_data_log_force[8299] <= 1'h0;
      write_enable_data_log_force[8300] <= 1'h0;
      write_enable_data_log_force[8301] <= 1'h0;
      write_enable_data_log_force[8302] <= 1'h0;
      write_enable_data_log_force[8303] <= 1'h0;
      write_enable_data_log_force[8304] <= 1'h0;
      write_enable_data_log_force[8305] <= 1'h0;
      write_enable_data_log_force[8306] <= 1'h0;
      write_enable_data_log_force[8307] <= 1'h0;
      write_enable_data_log_force[8308] <= 1'h0;
      write_enable_data_log_force[8309] <= 1'h0;
      write_enable_data_log_force[8310] <= 1'h0;
      write_enable_data_log_force[8311] <= 1'h0;
      write_enable_data_log_force[8312] <= 1'h0;
      write_enable_data_log_force[8313] <= 1'h0;
      write_enable_data_log_force[8314] <= 1'h0;
      write_enable_data_log_force[8315] <= 1'h0;
      write_enable_data_log_force[8316] <= 1'h0;
      write_enable_data_log_force[8317] <= 1'h0;
      write_enable_data_log_force[8318] <= 1'h0;
      write_enable_data_log_force[8319] <= 1'h0;

      // Input data for write_done_data_log
      write_done_data_log_force[   0] <= 1'h0;
      write_done_data_log_force[   1] <= 1'h0;
      write_done_data_log_force[   2] <= 1'h0;
      write_done_data_log_force[   3] <= 1'h0;
      write_done_data_log_force[   4] <= 1'h0;
      write_done_data_log_force[   5] <= 1'h0;
      write_done_data_log_force[   6] <= 1'h0;
      write_done_data_log_force[   7] <= 1'h0;
      write_done_data_log_force[   8] <= 1'h0;
      write_done_data_log_force[   9] <= 1'h0;
      write_done_data_log_force[  10] <= 1'h0;
      write_done_data_log_force[  11] <= 1'h0;
      write_done_data_log_force[  12] <= 1'h0;
      write_done_data_log_force[  13] <= 1'h0;
      write_done_data_log_force[  14] <= 1'h0;
      write_done_data_log_force[  15] <= 1'h0;
      write_done_data_log_force[  16] <= 1'h0;
      write_done_data_log_force[  17] <= 1'h0;
      write_done_data_log_force[  18] <= 1'h0;
      write_done_data_log_force[  19] <= 1'h0;
      write_done_data_log_force[  20] <= 1'h0;
      write_done_data_log_force[  21] <= 1'h0;
      write_done_data_log_force[  22] <= 1'h0;
      write_done_data_log_force[  23] <= 1'h0;
      write_done_data_log_force[  24] <= 1'h0;
      write_done_data_log_force[  25] <= 1'h0;
      write_done_data_log_force[  26] <= 1'h0;
      write_done_data_log_force[  27] <= 1'h0;
      write_done_data_log_force[  28] <= 1'h0;
      write_done_data_log_force[  29] <= 1'h0;
      write_done_data_log_force[  30] <= 1'h0;
      write_done_data_log_force[  31] <= 1'h0;
      write_done_data_log_force[  32] <= 1'h0;
      write_done_data_log_force[  33] <= 1'h0;
      write_done_data_log_force[  34] <= 1'h0;
      write_done_data_log_force[  35] <= 1'h0;
      write_done_data_log_force[  36] <= 1'h0;
      write_done_data_log_force[  37] <= 1'h0;
      write_done_data_log_force[  38] <= 1'h0;
      write_done_data_log_force[  39] <= 1'h0;
      write_done_data_log_force[  40] <= 1'h0;
      write_done_data_log_force[  41] <= 1'h0;
      write_done_data_log_force[  42] <= 1'h0;
      write_done_data_log_force[  43] <= 1'h0;
      write_done_data_log_force[  44] <= 1'h0;
      write_done_data_log_force[  45] <= 1'h0;
      write_done_data_log_force[  46] <= 1'h0;
      write_done_data_log_force[  47] <= 1'h0;
      write_done_data_log_force[  48] <= 1'h0;
      write_done_data_log_force[  49] <= 1'h0;
      write_done_data_log_force[  50] <= 1'h0;
      write_done_data_log_force[  51] <= 1'h0;
      write_done_data_log_force[  52] <= 1'h0;
      write_done_data_log_force[  53] <= 1'h0;
      write_done_data_log_force[  54] <= 1'h0;
      write_done_data_log_force[  55] <= 1'h0;
      write_done_data_log_force[  56] <= 1'h0;
      write_done_data_log_force[  57] <= 1'h0;
      write_done_data_log_force[  58] <= 1'h0;
      write_done_data_log_force[  59] <= 1'h0;
      write_done_data_log_force[  60] <= 1'h0;
      write_done_data_log_force[  61] <= 1'h0;
      write_done_data_log_force[  62] <= 1'h0;
      write_done_data_log_force[  63] <= 1'h0;
      write_done_data_log_force[  64] <= 1'h1;
      write_done_data_log_force[  65] <= 1'h0;
      write_done_data_log_force[  66] <= 1'h0;
      write_done_data_log_force[  67] <= 1'h0;
      write_done_data_log_force[  68] <= 1'h0;
      write_done_data_log_force[  69] <= 1'h0;
      write_done_data_log_force[  70] <= 1'h0;
      write_done_data_log_force[  71] <= 1'h0;
      write_done_data_log_force[  72] <= 1'h0;
      write_done_data_log_force[  73] <= 1'h0;
      write_done_data_log_force[  74] <= 1'h0;
      write_done_data_log_force[  75] <= 1'h0;
      write_done_data_log_force[  76] <= 1'h0;
      write_done_data_log_force[  77] <= 1'h0;
      write_done_data_log_force[  78] <= 1'h0;
      write_done_data_log_force[  79] <= 1'h0;
      write_done_data_log_force[  80] <= 1'h0;
      write_done_data_log_force[  81] <= 1'h0;
      write_done_data_log_force[  82] <= 1'h0;
      write_done_data_log_force[  83] <= 1'h0;
      write_done_data_log_force[  84] <= 1'h0;
      write_done_data_log_force[  85] <= 1'h0;
      write_done_data_log_force[  86] <= 1'h0;
      write_done_data_log_force[  87] <= 1'h0;
      write_done_data_log_force[  88] <= 1'h0;
      write_done_data_log_force[  89] <= 1'h0;
      write_done_data_log_force[  90] <= 1'h0;
      write_done_data_log_force[  91] <= 1'h0;
      write_done_data_log_force[  92] <= 1'h0;
      write_done_data_log_force[  93] <= 1'h0;
      write_done_data_log_force[  94] <= 1'h0;
      write_done_data_log_force[  95] <= 1'h0;
      write_done_data_log_force[  96] <= 1'h0;
      write_done_data_log_force[  97] <= 1'h0;
      write_done_data_log_force[  98] <= 1'h0;
      write_done_data_log_force[  99] <= 1'h0;
      write_done_data_log_force[ 100] <= 1'h0;
      write_done_data_log_force[ 101] <= 1'h0;
      write_done_data_log_force[ 102] <= 1'h0;
      write_done_data_log_force[ 103] <= 1'h0;
      write_done_data_log_force[ 104] <= 1'h0;
      write_done_data_log_force[ 105] <= 1'h0;
      write_done_data_log_force[ 106] <= 1'h0;
      write_done_data_log_force[ 107] <= 1'h0;
      write_done_data_log_force[ 108] <= 1'h0;
      write_done_data_log_force[ 109] <= 1'h0;
      write_done_data_log_force[ 110] <= 1'h0;
      write_done_data_log_force[ 111] <= 1'h0;
      write_done_data_log_force[ 112] <= 1'h0;
      write_done_data_log_force[ 113] <= 1'h0;
      write_done_data_log_force[ 114] <= 1'h0;
      write_done_data_log_force[ 115] <= 1'h0;
      write_done_data_log_force[ 116] <= 1'h0;
      write_done_data_log_force[ 117] <= 1'h0;
      write_done_data_log_force[ 118] <= 1'h0;
      write_done_data_log_force[ 119] <= 1'h0;
      write_done_data_log_force[ 120] <= 1'h0;
      write_done_data_log_force[ 121] <= 1'h0;
      write_done_data_log_force[ 122] <= 1'h0;
      write_done_data_log_force[ 123] <= 1'h0;
      write_done_data_log_force[ 124] <= 1'h0;
      write_done_data_log_force[ 125] <= 1'h0;
      write_done_data_log_force[ 126] <= 1'h0;
      write_done_data_log_force[ 127] <= 1'h0;
      write_done_data_log_force[ 128] <= 1'h0;
      write_done_data_log_force[ 129] <= 1'h0;
      write_done_data_log_force[ 130] <= 1'h0;
      write_done_data_log_force[ 131] <= 1'h0;
      write_done_data_log_force[ 132] <= 1'h0;
      write_done_data_log_force[ 133] <= 1'h0;
      write_done_data_log_force[ 134] <= 1'h0;
      write_done_data_log_force[ 135] <= 1'h0;
      write_done_data_log_force[ 136] <= 1'h0;
      write_done_data_log_force[ 137] <= 1'h0;
      write_done_data_log_force[ 138] <= 1'h0;
      write_done_data_log_force[ 139] <= 1'h0;
      write_done_data_log_force[ 140] <= 1'h0;
      write_done_data_log_force[ 141] <= 1'h0;
      write_done_data_log_force[ 142] <= 1'h0;
      write_done_data_log_force[ 143] <= 1'h0;
      write_done_data_log_force[ 144] <= 1'h0;
      write_done_data_log_force[ 145] <= 1'h0;
      write_done_data_log_force[ 146] <= 1'h0;
      write_done_data_log_force[ 147] <= 1'h0;
      write_done_data_log_force[ 148] <= 1'h0;
      write_done_data_log_force[ 149] <= 1'h0;
      write_done_data_log_force[ 150] <= 1'h0;
      write_done_data_log_force[ 151] <= 1'h0;
      write_done_data_log_force[ 152] <= 1'h0;
      write_done_data_log_force[ 153] <= 1'h0;
      write_done_data_log_force[ 154] <= 1'h0;
      write_done_data_log_force[ 155] <= 1'h0;
      write_done_data_log_force[ 156] <= 1'h0;
      write_done_data_log_force[ 157] <= 1'h0;
      write_done_data_log_force[ 158] <= 1'h0;
      write_done_data_log_force[ 159] <= 1'h0;
      write_done_data_log_force[ 160] <= 1'h0;
      write_done_data_log_force[ 161] <= 1'h0;
      write_done_data_log_force[ 162] <= 1'h0;
      write_done_data_log_force[ 163] <= 1'h0;
      write_done_data_log_force[ 164] <= 1'h0;
      write_done_data_log_force[ 165] <= 1'h0;
      write_done_data_log_force[ 166] <= 1'h0;
      write_done_data_log_force[ 167] <= 1'h0;
      write_done_data_log_force[ 168] <= 1'h0;
      write_done_data_log_force[ 169] <= 1'h0;
      write_done_data_log_force[ 170] <= 1'h0;
      write_done_data_log_force[ 171] <= 1'h0;
      write_done_data_log_force[ 172] <= 1'h0;
      write_done_data_log_force[ 173] <= 1'h0;
      write_done_data_log_force[ 174] <= 1'h0;
      write_done_data_log_force[ 175] <= 1'h0;
      write_done_data_log_force[ 176] <= 1'h0;
      write_done_data_log_force[ 177] <= 1'h0;
      write_done_data_log_force[ 178] <= 1'h0;
      write_done_data_log_force[ 179] <= 1'h0;
      write_done_data_log_force[ 180] <= 1'h0;
      write_done_data_log_force[ 181] <= 1'h0;
      write_done_data_log_force[ 182] <= 1'h0;
      write_done_data_log_force[ 183] <= 1'h0;
      write_done_data_log_force[ 184] <= 1'h0;
      write_done_data_log_force[ 185] <= 1'h0;
      write_done_data_log_force[ 186] <= 1'h0;
      write_done_data_log_force[ 187] <= 1'h0;
      write_done_data_log_force[ 188] <= 1'h0;
      write_done_data_log_force[ 189] <= 1'h0;
      write_done_data_log_force[ 190] <= 1'h0;
      write_done_data_log_force[ 191] <= 1'h0;
      write_done_data_log_force[ 192] <= 1'h0;
      write_done_data_log_force[ 193] <= 1'h0;
      write_done_data_log_force[ 194] <= 1'h0;
      write_done_data_log_force[ 195] <= 1'h0;
      write_done_data_log_force[ 196] <= 1'h0;
      write_done_data_log_force[ 197] <= 1'h0;
      write_done_data_log_force[ 198] <= 1'h0;
      write_done_data_log_force[ 199] <= 1'h0;
      write_done_data_log_force[ 200] <= 1'h0;
      write_done_data_log_force[ 201] <= 1'h0;
      write_done_data_log_force[ 202] <= 1'h0;
      write_done_data_log_force[ 203] <= 1'h0;
      write_done_data_log_force[ 204] <= 1'h0;
      write_done_data_log_force[ 205] <= 1'h0;
      write_done_data_log_force[ 206] <= 1'h0;
      write_done_data_log_force[ 207] <= 1'h0;
      write_done_data_log_force[ 208] <= 1'h0;
      write_done_data_log_force[ 209] <= 1'h0;
      write_done_data_log_force[ 210] <= 1'h0;
      write_done_data_log_force[ 211] <= 1'h0;
      write_done_data_log_force[ 212] <= 1'h0;
      write_done_data_log_force[ 213] <= 1'h0;
      write_done_data_log_force[ 214] <= 1'h0;
      write_done_data_log_force[ 215] <= 1'h0;
      write_done_data_log_force[ 216] <= 1'h0;
      write_done_data_log_force[ 217] <= 1'h0;
      write_done_data_log_force[ 218] <= 1'h0;
      write_done_data_log_force[ 219] <= 1'h0;
      write_done_data_log_force[ 220] <= 1'h0;
      write_done_data_log_force[ 221] <= 1'h0;
      write_done_data_log_force[ 222] <= 1'h0;
      write_done_data_log_force[ 223] <= 1'h0;
      write_done_data_log_force[ 224] <= 1'h0;
      write_done_data_log_force[ 225] <= 1'h0;
      write_done_data_log_force[ 226] <= 1'h0;
      write_done_data_log_force[ 227] <= 1'h0;
      write_done_data_log_force[ 228] <= 1'h0;
      write_done_data_log_force[ 229] <= 1'h0;
      write_done_data_log_force[ 230] <= 1'h0;
      write_done_data_log_force[ 231] <= 1'h0;
      write_done_data_log_force[ 232] <= 1'h0;
      write_done_data_log_force[ 233] <= 1'h0;
      write_done_data_log_force[ 234] <= 1'h0;
      write_done_data_log_force[ 235] <= 1'h0;
      write_done_data_log_force[ 236] <= 1'h0;
      write_done_data_log_force[ 237] <= 1'h0;
      write_done_data_log_force[ 238] <= 1'h0;
      write_done_data_log_force[ 239] <= 1'h0;
      write_done_data_log_force[ 240] <= 1'h0;
      write_done_data_log_force[ 241] <= 1'h0;
      write_done_data_log_force[ 242] <= 1'h0;
      write_done_data_log_force[ 243] <= 1'h0;
      write_done_data_log_force[ 244] <= 1'h0;
      write_done_data_log_force[ 245] <= 1'h0;
      write_done_data_log_force[ 246] <= 1'h0;
      write_done_data_log_force[ 247] <= 1'h0;
      write_done_data_log_force[ 248] <= 1'h0;
      write_done_data_log_force[ 249] <= 1'h0;
      write_done_data_log_force[ 250] <= 1'h0;
      write_done_data_log_force[ 251] <= 1'h0;
      write_done_data_log_force[ 252] <= 1'h0;
      write_done_data_log_force[ 253] <= 1'h0;
      write_done_data_log_force[ 254] <= 1'h0;
      write_done_data_log_force[ 255] <= 1'h0;
      write_done_data_log_force[ 256] <= 1'h0;
      write_done_data_log_force[ 257] <= 1'h0;
      write_done_data_log_force[ 258] <= 1'h0;
      write_done_data_log_force[ 259] <= 1'h0;
      write_done_data_log_force[ 260] <= 1'h0;
      write_done_data_log_force[ 261] <= 1'h0;
      write_done_data_log_force[ 262] <= 1'h0;
      write_done_data_log_force[ 263] <= 1'h0;
      write_done_data_log_force[ 264] <= 1'h0;
      write_done_data_log_force[ 265] <= 1'h0;
      write_done_data_log_force[ 266] <= 1'h0;
      write_done_data_log_force[ 267] <= 1'h0;
      write_done_data_log_force[ 268] <= 1'h0;
      write_done_data_log_force[ 269] <= 1'h0;
      write_done_data_log_force[ 270] <= 1'h0;
      write_done_data_log_force[ 271] <= 1'h0;
      write_done_data_log_force[ 272] <= 1'h0;
      write_done_data_log_force[ 273] <= 1'h0;
      write_done_data_log_force[ 274] <= 1'h0;
      write_done_data_log_force[ 275] <= 1'h0;
      write_done_data_log_force[ 276] <= 1'h0;
      write_done_data_log_force[ 277] <= 1'h0;
      write_done_data_log_force[ 278] <= 1'h0;
      write_done_data_log_force[ 279] <= 1'h0;
      write_done_data_log_force[ 280] <= 1'h0;
      write_done_data_log_force[ 281] <= 1'h0;
      write_done_data_log_force[ 282] <= 1'h0;
      write_done_data_log_force[ 283] <= 1'h0;
      write_done_data_log_force[ 284] <= 1'h0;
      write_done_data_log_force[ 285] <= 1'h0;
      write_done_data_log_force[ 286] <= 1'h0;
      write_done_data_log_force[ 287] <= 1'h0;
      write_done_data_log_force[ 288] <= 1'h0;
      write_done_data_log_force[ 289] <= 1'h0;
      write_done_data_log_force[ 290] <= 1'h0;
      write_done_data_log_force[ 291] <= 1'h0;
      write_done_data_log_force[ 292] <= 1'h0;
      write_done_data_log_force[ 293] <= 1'h0;
      write_done_data_log_force[ 294] <= 1'h0;
      write_done_data_log_force[ 295] <= 1'h0;
      write_done_data_log_force[ 296] <= 1'h0;
      write_done_data_log_force[ 297] <= 1'h0;
      write_done_data_log_force[ 298] <= 1'h0;
      write_done_data_log_force[ 299] <= 1'h0;
      write_done_data_log_force[ 300] <= 1'h0;
      write_done_data_log_force[ 301] <= 1'h0;
      write_done_data_log_force[ 302] <= 1'h0;
      write_done_data_log_force[ 303] <= 1'h0;
      write_done_data_log_force[ 304] <= 1'h0;
      write_done_data_log_force[ 305] <= 1'h0;
      write_done_data_log_force[ 306] <= 1'h0;
      write_done_data_log_force[ 307] <= 1'h0;
      write_done_data_log_force[ 308] <= 1'h0;
      write_done_data_log_force[ 309] <= 1'h0;
      write_done_data_log_force[ 310] <= 1'h0;
      write_done_data_log_force[ 311] <= 1'h0;
      write_done_data_log_force[ 312] <= 1'h0;
      write_done_data_log_force[ 313] <= 1'h0;
      write_done_data_log_force[ 314] <= 1'h0;
      write_done_data_log_force[ 315] <= 1'h0;
      write_done_data_log_force[ 316] <= 1'h0;
      write_done_data_log_force[ 317] <= 1'h0;
      write_done_data_log_force[ 318] <= 1'h0;
      write_done_data_log_force[ 319] <= 1'h0;
      write_done_data_log_force[ 320] <= 1'h0;
      write_done_data_log_force[ 321] <= 1'h0;
      write_done_data_log_force[ 322] <= 1'h0;
      write_done_data_log_force[ 323] <= 1'h0;
      write_done_data_log_force[ 324] <= 1'h0;
      write_done_data_log_force[ 325] <= 1'h0;
      write_done_data_log_force[ 326] <= 1'h0;
      write_done_data_log_force[ 327] <= 1'h0;
      write_done_data_log_force[ 328] <= 1'h0;
      write_done_data_log_force[ 329] <= 1'h0;
      write_done_data_log_force[ 330] <= 1'h0;
      write_done_data_log_force[ 331] <= 1'h0;
      write_done_data_log_force[ 332] <= 1'h0;
      write_done_data_log_force[ 333] <= 1'h0;
      write_done_data_log_force[ 334] <= 1'h0;
      write_done_data_log_force[ 335] <= 1'h0;
      write_done_data_log_force[ 336] <= 1'h0;
      write_done_data_log_force[ 337] <= 1'h0;
      write_done_data_log_force[ 338] <= 1'h0;
      write_done_data_log_force[ 339] <= 1'h0;
      write_done_data_log_force[ 340] <= 1'h0;
      write_done_data_log_force[ 341] <= 1'h0;
      write_done_data_log_force[ 342] <= 1'h0;
      write_done_data_log_force[ 343] <= 1'h0;
      write_done_data_log_force[ 344] <= 1'h0;
      write_done_data_log_force[ 345] <= 1'h0;
      write_done_data_log_force[ 346] <= 1'h0;
      write_done_data_log_force[ 347] <= 1'h0;
      write_done_data_log_force[ 348] <= 1'h0;
      write_done_data_log_force[ 349] <= 1'h0;
      write_done_data_log_force[ 350] <= 1'h0;
      write_done_data_log_force[ 351] <= 1'h0;
      write_done_data_log_force[ 352] <= 1'h0;
      write_done_data_log_force[ 353] <= 1'h0;
      write_done_data_log_force[ 354] <= 1'h0;
      write_done_data_log_force[ 355] <= 1'h0;
      write_done_data_log_force[ 356] <= 1'h0;
      write_done_data_log_force[ 357] <= 1'h0;
      write_done_data_log_force[ 358] <= 1'h0;
      write_done_data_log_force[ 359] <= 1'h0;
      write_done_data_log_force[ 360] <= 1'h0;
      write_done_data_log_force[ 361] <= 1'h0;
      write_done_data_log_force[ 362] <= 1'h0;
      write_done_data_log_force[ 363] <= 1'h0;
      write_done_data_log_force[ 364] <= 1'h0;
      write_done_data_log_force[ 365] <= 1'h0;
      write_done_data_log_force[ 366] <= 1'h0;
      write_done_data_log_force[ 367] <= 1'h0;
      write_done_data_log_force[ 368] <= 1'h0;
      write_done_data_log_force[ 369] <= 1'h0;
      write_done_data_log_force[ 370] <= 1'h0;
      write_done_data_log_force[ 371] <= 1'h0;
      write_done_data_log_force[ 372] <= 1'h0;
      write_done_data_log_force[ 373] <= 1'h0;
      write_done_data_log_force[ 374] <= 1'h0;
      write_done_data_log_force[ 375] <= 1'h0;
      write_done_data_log_force[ 376] <= 1'h0;
      write_done_data_log_force[ 377] <= 1'h0;
      write_done_data_log_force[ 378] <= 1'h0;
      write_done_data_log_force[ 379] <= 1'h0;
      write_done_data_log_force[ 380] <= 1'h0;
      write_done_data_log_force[ 381] <= 1'h0;
      write_done_data_log_force[ 382] <= 1'h0;
      write_done_data_log_force[ 383] <= 1'h0;
      write_done_data_log_force[ 384] <= 1'h0;
      write_done_data_log_force[ 385] <= 1'h0;
      write_done_data_log_force[ 386] <= 1'h0;
      write_done_data_log_force[ 387] <= 1'h0;
      write_done_data_log_force[ 388] <= 1'h0;
      write_done_data_log_force[ 389] <= 1'h0;
      write_done_data_log_force[ 390] <= 1'h0;
      write_done_data_log_force[ 391] <= 1'h0;
      write_done_data_log_force[ 392] <= 1'h0;
      write_done_data_log_force[ 393] <= 1'h0;
      write_done_data_log_force[ 394] <= 1'h0;
      write_done_data_log_force[ 395] <= 1'h0;
      write_done_data_log_force[ 396] <= 1'h0;
      write_done_data_log_force[ 397] <= 1'h0;
      write_done_data_log_force[ 398] <= 1'h0;
      write_done_data_log_force[ 399] <= 1'h0;
      write_done_data_log_force[ 400] <= 1'h0;
      write_done_data_log_force[ 401] <= 1'h0;
      write_done_data_log_force[ 402] <= 1'h0;
      write_done_data_log_force[ 403] <= 1'h0;
      write_done_data_log_force[ 404] <= 1'h0;
      write_done_data_log_force[ 405] <= 1'h0;
      write_done_data_log_force[ 406] <= 1'h0;
      write_done_data_log_force[ 407] <= 1'h0;
      write_done_data_log_force[ 408] <= 1'h0;
      write_done_data_log_force[ 409] <= 1'h0;
      write_done_data_log_force[ 410] <= 1'h0;
      write_done_data_log_force[ 411] <= 1'h0;
      write_done_data_log_force[ 412] <= 1'h0;
      write_done_data_log_force[ 413] <= 1'h0;
      write_done_data_log_force[ 414] <= 1'h0;
      write_done_data_log_force[ 415] <= 1'h0;
      write_done_data_log_force[ 416] <= 1'h0;
      write_done_data_log_force[ 417] <= 1'h0;
      write_done_data_log_force[ 418] <= 1'h0;
      write_done_data_log_force[ 419] <= 1'h0;
      write_done_data_log_force[ 420] <= 1'h0;
      write_done_data_log_force[ 421] <= 1'h0;
      write_done_data_log_force[ 422] <= 1'h0;
      write_done_data_log_force[ 423] <= 1'h0;
      write_done_data_log_force[ 424] <= 1'h0;
      write_done_data_log_force[ 425] <= 1'h0;
      write_done_data_log_force[ 426] <= 1'h0;
      write_done_data_log_force[ 427] <= 1'h0;
      write_done_data_log_force[ 428] <= 1'h0;
      write_done_data_log_force[ 429] <= 1'h0;
      write_done_data_log_force[ 430] <= 1'h0;
      write_done_data_log_force[ 431] <= 1'h0;
      write_done_data_log_force[ 432] <= 1'h0;
      write_done_data_log_force[ 433] <= 1'h0;
      write_done_data_log_force[ 434] <= 1'h0;
      write_done_data_log_force[ 435] <= 1'h0;
      write_done_data_log_force[ 436] <= 1'h0;
      write_done_data_log_force[ 437] <= 1'h0;
      write_done_data_log_force[ 438] <= 1'h0;
      write_done_data_log_force[ 439] <= 1'h0;
      write_done_data_log_force[ 440] <= 1'h0;
      write_done_data_log_force[ 441] <= 1'h0;
      write_done_data_log_force[ 442] <= 1'h0;
      write_done_data_log_force[ 443] <= 1'h0;
      write_done_data_log_force[ 444] <= 1'h0;
      write_done_data_log_force[ 445] <= 1'h0;
      write_done_data_log_force[ 446] <= 1'h0;
      write_done_data_log_force[ 447] <= 1'h0;
      write_done_data_log_force[ 448] <= 1'h0;
      write_done_data_log_force[ 449] <= 1'h0;
      write_done_data_log_force[ 450] <= 1'h0;
      write_done_data_log_force[ 451] <= 1'h0;
      write_done_data_log_force[ 452] <= 1'h0;
      write_done_data_log_force[ 453] <= 1'h0;
      write_done_data_log_force[ 454] <= 1'h0;
      write_done_data_log_force[ 455] <= 1'h0;
      write_done_data_log_force[ 456] <= 1'h0;
      write_done_data_log_force[ 457] <= 1'h0;
      write_done_data_log_force[ 458] <= 1'h0;
      write_done_data_log_force[ 459] <= 1'h0;
      write_done_data_log_force[ 460] <= 1'h0;
      write_done_data_log_force[ 461] <= 1'h0;
      write_done_data_log_force[ 462] <= 1'h0;
      write_done_data_log_force[ 463] <= 1'h0;
      write_done_data_log_force[ 464] <= 1'h0;
      write_done_data_log_force[ 465] <= 1'h0;
      write_done_data_log_force[ 466] <= 1'h0;
      write_done_data_log_force[ 467] <= 1'h0;
      write_done_data_log_force[ 468] <= 1'h0;
      write_done_data_log_force[ 469] <= 1'h0;
      write_done_data_log_force[ 470] <= 1'h0;
      write_done_data_log_force[ 471] <= 1'h0;
      write_done_data_log_force[ 472] <= 1'h0;
      write_done_data_log_force[ 473] <= 1'h0;
      write_done_data_log_force[ 474] <= 1'h0;
      write_done_data_log_force[ 475] <= 1'h0;
      write_done_data_log_force[ 476] <= 1'h0;
      write_done_data_log_force[ 477] <= 1'h0;
      write_done_data_log_force[ 478] <= 1'h0;
      write_done_data_log_force[ 479] <= 1'h0;
      write_done_data_log_force[ 480] <= 1'h0;
      write_done_data_log_force[ 481] <= 1'h0;
      write_done_data_log_force[ 482] <= 1'h0;
      write_done_data_log_force[ 483] <= 1'h0;
      write_done_data_log_force[ 484] <= 1'h0;
      write_done_data_log_force[ 485] <= 1'h0;
      write_done_data_log_force[ 486] <= 1'h0;
      write_done_data_log_force[ 487] <= 1'h0;
      write_done_data_log_force[ 488] <= 1'h0;
      write_done_data_log_force[ 489] <= 1'h0;
      write_done_data_log_force[ 490] <= 1'h0;
      write_done_data_log_force[ 491] <= 1'h0;
      write_done_data_log_force[ 492] <= 1'h0;
      write_done_data_log_force[ 493] <= 1'h0;
      write_done_data_log_force[ 494] <= 1'h0;
      write_done_data_log_force[ 495] <= 1'h0;
      write_done_data_log_force[ 496] <= 1'h0;
      write_done_data_log_force[ 497] <= 1'h0;
      write_done_data_log_force[ 498] <= 1'h0;
      write_done_data_log_force[ 499] <= 1'h0;
      write_done_data_log_force[ 500] <= 1'h0;
      write_done_data_log_force[ 501] <= 1'h0;
      write_done_data_log_force[ 502] <= 1'h0;
      write_done_data_log_force[ 503] <= 1'h0;
      write_done_data_log_force[ 504] <= 1'h0;
      write_done_data_log_force[ 505] <= 1'h0;
      write_done_data_log_force[ 506] <= 1'h0;
      write_done_data_log_force[ 507] <= 1'h0;
      write_done_data_log_force[ 508] <= 1'h0;
      write_done_data_log_force[ 509] <= 1'h0;
      write_done_data_log_force[ 510] <= 1'h0;
      write_done_data_log_force[ 511] <= 1'h0;
      write_done_data_log_force[ 512] <= 1'h0;
      write_done_data_log_force[ 513] <= 1'h0;
      write_done_data_log_force[ 514] <= 1'h0;
      write_done_data_log_force[ 515] <= 1'h0;
      write_done_data_log_force[ 516] <= 1'h0;
      write_done_data_log_force[ 517] <= 1'h0;
      write_done_data_log_force[ 518] <= 1'h0;
      write_done_data_log_force[ 519] <= 1'h0;
      write_done_data_log_force[ 520] <= 1'h0;
      write_done_data_log_force[ 521] <= 1'h0;
      write_done_data_log_force[ 522] <= 1'h0;
      write_done_data_log_force[ 523] <= 1'h0;
      write_done_data_log_force[ 524] <= 1'h0;
      write_done_data_log_force[ 525] <= 1'h0;
      write_done_data_log_force[ 526] <= 1'h0;
      write_done_data_log_force[ 527] <= 1'h0;
      write_done_data_log_force[ 528] <= 1'h0;
      write_done_data_log_force[ 529] <= 1'h0;
      write_done_data_log_force[ 530] <= 1'h0;
      write_done_data_log_force[ 531] <= 1'h0;
      write_done_data_log_force[ 532] <= 1'h0;
      write_done_data_log_force[ 533] <= 1'h0;
      write_done_data_log_force[ 534] <= 1'h0;
      write_done_data_log_force[ 535] <= 1'h0;
      write_done_data_log_force[ 536] <= 1'h0;
      write_done_data_log_force[ 537] <= 1'h0;
      write_done_data_log_force[ 538] <= 1'h0;
      write_done_data_log_force[ 539] <= 1'h0;
      write_done_data_log_force[ 540] <= 1'h0;
      write_done_data_log_force[ 541] <= 1'h0;
      write_done_data_log_force[ 542] <= 1'h0;
      write_done_data_log_force[ 543] <= 1'h0;
      write_done_data_log_force[ 544] <= 1'h0;
      write_done_data_log_force[ 545] <= 1'h0;
      write_done_data_log_force[ 546] <= 1'h0;
      write_done_data_log_force[ 547] <= 1'h0;
      write_done_data_log_force[ 548] <= 1'h0;
      write_done_data_log_force[ 549] <= 1'h0;
      write_done_data_log_force[ 550] <= 1'h0;
      write_done_data_log_force[ 551] <= 1'h0;
      write_done_data_log_force[ 552] <= 1'h0;
      write_done_data_log_force[ 553] <= 1'h0;
      write_done_data_log_force[ 554] <= 1'h0;
      write_done_data_log_force[ 555] <= 1'h0;
      write_done_data_log_force[ 556] <= 1'h0;
      write_done_data_log_force[ 557] <= 1'h0;
      write_done_data_log_force[ 558] <= 1'h0;
      write_done_data_log_force[ 559] <= 1'h0;
      write_done_data_log_force[ 560] <= 1'h0;
      write_done_data_log_force[ 561] <= 1'h0;
      write_done_data_log_force[ 562] <= 1'h0;
      write_done_data_log_force[ 563] <= 1'h0;
      write_done_data_log_force[ 564] <= 1'h0;
      write_done_data_log_force[ 565] <= 1'h0;
      write_done_data_log_force[ 566] <= 1'h0;
      write_done_data_log_force[ 567] <= 1'h0;
      write_done_data_log_force[ 568] <= 1'h0;
      write_done_data_log_force[ 569] <= 1'h0;
      write_done_data_log_force[ 570] <= 1'h0;
      write_done_data_log_force[ 571] <= 1'h0;
      write_done_data_log_force[ 572] <= 1'h0;
      write_done_data_log_force[ 573] <= 1'h0;
      write_done_data_log_force[ 574] <= 1'h0;
      write_done_data_log_force[ 575] <= 1'h0;
      write_done_data_log_force[ 576] <= 1'h0;
      write_done_data_log_force[ 577] <= 1'h0;
      write_done_data_log_force[ 578] <= 1'h0;
      write_done_data_log_force[ 579] <= 1'h0;
      write_done_data_log_force[ 580] <= 1'h0;
      write_done_data_log_force[ 581] <= 1'h0;
      write_done_data_log_force[ 582] <= 1'h0;
      write_done_data_log_force[ 583] <= 1'h0;
      write_done_data_log_force[ 584] <= 1'h0;
      write_done_data_log_force[ 585] <= 1'h0;
      write_done_data_log_force[ 586] <= 1'h0;
      write_done_data_log_force[ 587] <= 1'h0;
      write_done_data_log_force[ 588] <= 1'h0;
      write_done_data_log_force[ 589] <= 1'h0;
      write_done_data_log_force[ 590] <= 1'h0;
      write_done_data_log_force[ 591] <= 1'h0;
      write_done_data_log_force[ 592] <= 1'h0;
      write_done_data_log_force[ 593] <= 1'h0;
      write_done_data_log_force[ 594] <= 1'h0;
      write_done_data_log_force[ 595] <= 1'h0;
      write_done_data_log_force[ 596] <= 1'h0;
      write_done_data_log_force[ 597] <= 1'h0;
      write_done_data_log_force[ 598] <= 1'h0;
      write_done_data_log_force[ 599] <= 1'h0;
      write_done_data_log_force[ 600] <= 1'h0;
      write_done_data_log_force[ 601] <= 1'h0;
      write_done_data_log_force[ 602] <= 1'h0;
      write_done_data_log_force[ 603] <= 1'h0;
      write_done_data_log_force[ 604] <= 1'h0;
      write_done_data_log_force[ 605] <= 1'h0;
      write_done_data_log_force[ 606] <= 1'h0;
      write_done_data_log_force[ 607] <= 1'h0;
      write_done_data_log_force[ 608] <= 1'h0;
      write_done_data_log_force[ 609] <= 1'h0;
      write_done_data_log_force[ 610] <= 1'h0;
      write_done_data_log_force[ 611] <= 1'h0;
      write_done_data_log_force[ 612] <= 1'h0;
      write_done_data_log_force[ 613] <= 1'h0;
      write_done_data_log_force[ 614] <= 1'h0;
      write_done_data_log_force[ 615] <= 1'h0;
      write_done_data_log_force[ 616] <= 1'h0;
      write_done_data_log_force[ 617] <= 1'h0;
      write_done_data_log_force[ 618] <= 1'h0;
      write_done_data_log_force[ 619] <= 1'h0;
      write_done_data_log_force[ 620] <= 1'h0;
      write_done_data_log_force[ 621] <= 1'h0;
      write_done_data_log_force[ 622] <= 1'h0;
      write_done_data_log_force[ 623] <= 1'h0;
      write_done_data_log_force[ 624] <= 1'h0;
      write_done_data_log_force[ 625] <= 1'h0;
      write_done_data_log_force[ 626] <= 1'h0;
      write_done_data_log_force[ 627] <= 1'h0;
      write_done_data_log_force[ 628] <= 1'h0;
      write_done_data_log_force[ 629] <= 1'h0;
      write_done_data_log_force[ 630] <= 1'h0;
      write_done_data_log_force[ 631] <= 1'h0;
      write_done_data_log_force[ 632] <= 1'h0;
      write_done_data_log_force[ 633] <= 1'h0;
      write_done_data_log_force[ 634] <= 1'h0;
      write_done_data_log_force[ 635] <= 1'h0;
      write_done_data_log_force[ 636] <= 1'h0;
      write_done_data_log_force[ 637] <= 1'h0;
      write_done_data_log_force[ 638] <= 1'h0;
      write_done_data_log_force[ 639] <= 1'h0;
      write_done_data_log_force[ 640] <= 1'h0;
      write_done_data_log_force[ 641] <= 1'h0;
      write_done_data_log_force[ 642] <= 1'h0;
      write_done_data_log_force[ 643] <= 1'h0;
      write_done_data_log_force[ 644] <= 1'h0;
      write_done_data_log_force[ 645] <= 1'h0;
      write_done_data_log_force[ 646] <= 1'h0;
      write_done_data_log_force[ 647] <= 1'h0;
      write_done_data_log_force[ 648] <= 1'h0;
      write_done_data_log_force[ 649] <= 1'h0;
      write_done_data_log_force[ 650] <= 1'h0;
      write_done_data_log_force[ 651] <= 1'h0;
      write_done_data_log_force[ 652] <= 1'h0;
      write_done_data_log_force[ 653] <= 1'h0;
      write_done_data_log_force[ 654] <= 1'h0;
      write_done_data_log_force[ 655] <= 1'h0;
      write_done_data_log_force[ 656] <= 1'h0;
      write_done_data_log_force[ 657] <= 1'h0;
      write_done_data_log_force[ 658] <= 1'h0;
      write_done_data_log_force[ 659] <= 1'h0;
      write_done_data_log_force[ 660] <= 1'h0;
      write_done_data_log_force[ 661] <= 1'h0;
      write_done_data_log_force[ 662] <= 1'h0;
      write_done_data_log_force[ 663] <= 1'h0;
      write_done_data_log_force[ 664] <= 1'h0;
      write_done_data_log_force[ 665] <= 1'h0;
      write_done_data_log_force[ 666] <= 1'h0;
      write_done_data_log_force[ 667] <= 1'h0;
      write_done_data_log_force[ 668] <= 1'h0;
      write_done_data_log_force[ 669] <= 1'h0;
      write_done_data_log_force[ 670] <= 1'h0;
      write_done_data_log_force[ 671] <= 1'h0;
      write_done_data_log_force[ 672] <= 1'h0;
      write_done_data_log_force[ 673] <= 1'h0;
      write_done_data_log_force[ 674] <= 1'h0;
      write_done_data_log_force[ 675] <= 1'h0;
      write_done_data_log_force[ 676] <= 1'h0;
      write_done_data_log_force[ 677] <= 1'h0;
      write_done_data_log_force[ 678] <= 1'h0;
      write_done_data_log_force[ 679] <= 1'h0;
      write_done_data_log_force[ 680] <= 1'h0;
      write_done_data_log_force[ 681] <= 1'h0;
      write_done_data_log_force[ 682] <= 1'h0;
      write_done_data_log_force[ 683] <= 1'h0;
      write_done_data_log_force[ 684] <= 1'h0;
      write_done_data_log_force[ 685] <= 1'h0;
      write_done_data_log_force[ 686] <= 1'h0;
      write_done_data_log_force[ 687] <= 1'h0;
      write_done_data_log_force[ 688] <= 1'h0;
      write_done_data_log_force[ 689] <= 1'h0;
      write_done_data_log_force[ 690] <= 1'h0;
      write_done_data_log_force[ 691] <= 1'h0;
      write_done_data_log_force[ 692] <= 1'h0;
      write_done_data_log_force[ 693] <= 1'h0;
      write_done_data_log_force[ 694] <= 1'h0;
      write_done_data_log_force[ 695] <= 1'h0;
      write_done_data_log_force[ 696] <= 1'h0;
      write_done_data_log_force[ 697] <= 1'h0;
      write_done_data_log_force[ 698] <= 1'h0;
      write_done_data_log_force[ 699] <= 1'h0;
      write_done_data_log_force[ 700] <= 1'h0;
      write_done_data_log_force[ 701] <= 1'h0;
      write_done_data_log_force[ 702] <= 1'h0;
      write_done_data_log_force[ 703] <= 1'h0;
      write_done_data_log_force[ 704] <= 1'h0;
      write_done_data_log_force[ 705] <= 1'h0;
      write_done_data_log_force[ 706] <= 1'h0;
      write_done_data_log_force[ 707] <= 1'h0;
      write_done_data_log_force[ 708] <= 1'h0;
      write_done_data_log_force[ 709] <= 1'h0;
      write_done_data_log_force[ 710] <= 1'h0;
      write_done_data_log_force[ 711] <= 1'h0;
      write_done_data_log_force[ 712] <= 1'h0;
      write_done_data_log_force[ 713] <= 1'h0;
      write_done_data_log_force[ 714] <= 1'h0;
      write_done_data_log_force[ 715] <= 1'h0;
      write_done_data_log_force[ 716] <= 1'h0;
      write_done_data_log_force[ 717] <= 1'h0;
      write_done_data_log_force[ 718] <= 1'h0;
      write_done_data_log_force[ 719] <= 1'h0;
      write_done_data_log_force[ 720] <= 1'h0;
      write_done_data_log_force[ 721] <= 1'h0;
      write_done_data_log_force[ 722] <= 1'h0;
      write_done_data_log_force[ 723] <= 1'h0;
      write_done_data_log_force[ 724] <= 1'h0;
      write_done_data_log_force[ 725] <= 1'h0;
      write_done_data_log_force[ 726] <= 1'h0;
      write_done_data_log_force[ 727] <= 1'h0;
      write_done_data_log_force[ 728] <= 1'h0;
      write_done_data_log_force[ 729] <= 1'h0;
      write_done_data_log_force[ 730] <= 1'h0;
      write_done_data_log_force[ 731] <= 1'h0;
      write_done_data_log_force[ 732] <= 1'h0;
      write_done_data_log_force[ 733] <= 1'h0;
      write_done_data_log_force[ 734] <= 1'h0;
      write_done_data_log_force[ 735] <= 1'h0;
      write_done_data_log_force[ 736] <= 1'h0;
      write_done_data_log_force[ 737] <= 1'h0;
      write_done_data_log_force[ 738] <= 1'h0;
      write_done_data_log_force[ 739] <= 1'h0;
      write_done_data_log_force[ 740] <= 1'h0;
      write_done_data_log_force[ 741] <= 1'h0;
      write_done_data_log_force[ 742] <= 1'h0;
      write_done_data_log_force[ 743] <= 1'h0;
      write_done_data_log_force[ 744] <= 1'h0;
      write_done_data_log_force[ 745] <= 1'h0;
      write_done_data_log_force[ 746] <= 1'h0;
      write_done_data_log_force[ 747] <= 1'h0;
      write_done_data_log_force[ 748] <= 1'h0;
      write_done_data_log_force[ 749] <= 1'h0;
      write_done_data_log_force[ 750] <= 1'h0;
      write_done_data_log_force[ 751] <= 1'h0;
      write_done_data_log_force[ 752] <= 1'h0;
      write_done_data_log_force[ 753] <= 1'h0;
      write_done_data_log_force[ 754] <= 1'h0;
      write_done_data_log_force[ 755] <= 1'h0;
      write_done_data_log_force[ 756] <= 1'h0;
      write_done_data_log_force[ 757] <= 1'h0;
      write_done_data_log_force[ 758] <= 1'h0;
      write_done_data_log_force[ 759] <= 1'h0;
      write_done_data_log_force[ 760] <= 1'h0;
      write_done_data_log_force[ 761] <= 1'h0;
      write_done_data_log_force[ 762] <= 1'h0;
      write_done_data_log_force[ 763] <= 1'h0;
      write_done_data_log_force[ 764] <= 1'h0;
      write_done_data_log_force[ 765] <= 1'h0;
      write_done_data_log_force[ 766] <= 1'h0;
      write_done_data_log_force[ 767] <= 1'h0;
      write_done_data_log_force[ 768] <= 1'h0;
      write_done_data_log_force[ 769] <= 1'h0;
      write_done_data_log_force[ 770] <= 1'h0;
      write_done_data_log_force[ 771] <= 1'h0;
      write_done_data_log_force[ 772] <= 1'h0;
      write_done_data_log_force[ 773] <= 1'h0;
      write_done_data_log_force[ 774] <= 1'h0;
      write_done_data_log_force[ 775] <= 1'h0;
      write_done_data_log_force[ 776] <= 1'h0;
      write_done_data_log_force[ 777] <= 1'h0;
      write_done_data_log_force[ 778] <= 1'h0;
      write_done_data_log_force[ 779] <= 1'h0;
      write_done_data_log_force[ 780] <= 1'h0;
      write_done_data_log_force[ 781] <= 1'h0;
      write_done_data_log_force[ 782] <= 1'h0;
      write_done_data_log_force[ 783] <= 1'h0;
      write_done_data_log_force[ 784] <= 1'h0;
      write_done_data_log_force[ 785] <= 1'h0;
      write_done_data_log_force[ 786] <= 1'h0;
      write_done_data_log_force[ 787] <= 1'h0;
      write_done_data_log_force[ 788] <= 1'h0;
      write_done_data_log_force[ 789] <= 1'h0;
      write_done_data_log_force[ 790] <= 1'h0;
      write_done_data_log_force[ 791] <= 1'h0;
      write_done_data_log_force[ 792] <= 1'h0;
      write_done_data_log_force[ 793] <= 1'h0;
      write_done_data_log_force[ 794] <= 1'h0;
      write_done_data_log_force[ 795] <= 1'h0;
      write_done_data_log_force[ 796] <= 1'h0;
      write_done_data_log_force[ 797] <= 1'h0;
      write_done_data_log_force[ 798] <= 1'h0;
      write_done_data_log_force[ 799] <= 1'h0;
      write_done_data_log_force[ 800] <= 1'h0;
      write_done_data_log_force[ 801] <= 1'h0;
      write_done_data_log_force[ 802] <= 1'h0;
      write_done_data_log_force[ 803] <= 1'h0;
      write_done_data_log_force[ 804] <= 1'h0;
      write_done_data_log_force[ 805] <= 1'h0;
      write_done_data_log_force[ 806] <= 1'h0;
      write_done_data_log_force[ 807] <= 1'h0;
      write_done_data_log_force[ 808] <= 1'h0;
      write_done_data_log_force[ 809] <= 1'h0;
      write_done_data_log_force[ 810] <= 1'h0;
      write_done_data_log_force[ 811] <= 1'h0;
      write_done_data_log_force[ 812] <= 1'h0;
      write_done_data_log_force[ 813] <= 1'h0;
      write_done_data_log_force[ 814] <= 1'h0;
      write_done_data_log_force[ 815] <= 1'h0;
      write_done_data_log_force[ 816] <= 1'h0;
      write_done_data_log_force[ 817] <= 1'h0;
      write_done_data_log_force[ 818] <= 1'h0;
      write_done_data_log_force[ 819] <= 1'h0;
      write_done_data_log_force[ 820] <= 1'h0;
      write_done_data_log_force[ 821] <= 1'h0;
      write_done_data_log_force[ 822] <= 1'h0;
      write_done_data_log_force[ 823] <= 1'h0;
      write_done_data_log_force[ 824] <= 1'h0;
      write_done_data_log_force[ 825] <= 1'h0;
      write_done_data_log_force[ 826] <= 1'h0;
      write_done_data_log_force[ 827] <= 1'h0;
      write_done_data_log_force[ 828] <= 1'h0;
      write_done_data_log_force[ 829] <= 1'h0;
      write_done_data_log_force[ 830] <= 1'h0;
      write_done_data_log_force[ 831] <= 1'h0;
      write_done_data_log_force[ 832] <= 1'h0;
      write_done_data_log_force[ 833] <= 1'h0;
      write_done_data_log_force[ 834] <= 1'h0;
      write_done_data_log_force[ 835] <= 1'h0;
      write_done_data_log_force[ 836] <= 1'h0;
      write_done_data_log_force[ 837] <= 1'h0;
      write_done_data_log_force[ 838] <= 1'h0;
      write_done_data_log_force[ 839] <= 1'h0;
      write_done_data_log_force[ 840] <= 1'h0;
      write_done_data_log_force[ 841] <= 1'h0;
      write_done_data_log_force[ 842] <= 1'h0;
      write_done_data_log_force[ 843] <= 1'h0;
      write_done_data_log_force[ 844] <= 1'h0;
      write_done_data_log_force[ 845] <= 1'h0;
      write_done_data_log_force[ 846] <= 1'h0;
      write_done_data_log_force[ 847] <= 1'h0;
      write_done_data_log_force[ 848] <= 1'h0;
      write_done_data_log_force[ 849] <= 1'h0;
      write_done_data_log_force[ 850] <= 1'h0;
      write_done_data_log_force[ 851] <= 1'h0;
      write_done_data_log_force[ 852] <= 1'h0;
      write_done_data_log_force[ 853] <= 1'h0;
      write_done_data_log_force[ 854] <= 1'h0;
      write_done_data_log_force[ 855] <= 1'h0;
      write_done_data_log_force[ 856] <= 1'h0;
      write_done_data_log_force[ 857] <= 1'h0;
      write_done_data_log_force[ 858] <= 1'h0;
      write_done_data_log_force[ 859] <= 1'h0;
      write_done_data_log_force[ 860] <= 1'h0;
      write_done_data_log_force[ 861] <= 1'h0;
      write_done_data_log_force[ 862] <= 1'h0;
      write_done_data_log_force[ 863] <= 1'h0;
      write_done_data_log_force[ 864] <= 1'h0;
      write_done_data_log_force[ 865] <= 1'h0;
      write_done_data_log_force[ 866] <= 1'h0;
      write_done_data_log_force[ 867] <= 1'h0;
      write_done_data_log_force[ 868] <= 1'h0;
      write_done_data_log_force[ 869] <= 1'h0;
      write_done_data_log_force[ 870] <= 1'h0;
      write_done_data_log_force[ 871] <= 1'h0;
      write_done_data_log_force[ 872] <= 1'h0;
      write_done_data_log_force[ 873] <= 1'h0;
      write_done_data_log_force[ 874] <= 1'h0;
      write_done_data_log_force[ 875] <= 1'h0;
      write_done_data_log_force[ 876] <= 1'h0;
      write_done_data_log_force[ 877] <= 1'h0;
      write_done_data_log_force[ 878] <= 1'h0;
      write_done_data_log_force[ 879] <= 1'h0;
      write_done_data_log_force[ 880] <= 1'h0;
      write_done_data_log_force[ 881] <= 1'h0;
      write_done_data_log_force[ 882] <= 1'h0;
      write_done_data_log_force[ 883] <= 1'h0;
      write_done_data_log_force[ 884] <= 1'h0;
      write_done_data_log_force[ 885] <= 1'h0;
      write_done_data_log_force[ 886] <= 1'h0;
      write_done_data_log_force[ 887] <= 1'h0;
      write_done_data_log_force[ 888] <= 1'h0;
      write_done_data_log_force[ 889] <= 1'h0;
      write_done_data_log_force[ 890] <= 1'h0;
      write_done_data_log_force[ 891] <= 1'h0;
      write_done_data_log_force[ 892] <= 1'h0;
      write_done_data_log_force[ 893] <= 1'h0;
      write_done_data_log_force[ 894] <= 1'h0;
      write_done_data_log_force[ 895] <= 1'h0;
      write_done_data_log_force[ 896] <= 1'h0;
      write_done_data_log_force[ 897] <= 1'h0;
      write_done_data_log_force[ 898] <= 1'h0;
      write_done_data_log_force[ 899] <= 1'h0;
      write_done_data_log_force[ 900] <= 1'h0;
      write_done_data_log_force[ 901] <= 1'h0;
      write_done_data_log_force[ 902] <= 1'h0;
      write_done_data_log_force[ 903] <= 1'h0;
      write_done_data_log_force[ 904] <= 1'h0;
      write_done_data_log_force[ 905] <= 1'h0;
      write_done_data_log_force[ 906] <= 1'h0;
      write_done_data_log_force[ 907] <= 1'h0;
      write_done_data_log_force[ 908] <= 1'h0;
      write_done_data_log_force[ 909] <= 1'h0;
      write_done_data_log_force[ 910] <= 1'h0;
      write_done_data_log_force[ 911] <= 1'h0;
      write_done_data_log_force[ 912] <= 1'h0;
      write_done_data_log_force[ 913] <= 1'h0;
      write_done_data_log_force[ 914] <= 1'h0;
      write_done_data_log_force[ 915] <= 1'h0;
      write_done_data_log_force[ 916] <= 1'h0;
      write_done_data_log_force[ 917] <= 1'h0;
      write_done_data_log_force[ 918] <= 1'h0;
      write_done_data_log_force[ 919] <= 1'h0;
      write_done_data_log_force[ 920] <= 1'h0;
      write_done_data_log_force[ 921] <= 1'h0;
      write_done_data_log_force[ 922] <= 1'h0;
      write_done_data_log_force[ 923] <= 1'h0;
      write_done_data_log_force[ 924] <= 1'h0;
      write_done_data_log_force[ 925] <= 1'h0;
      write_done_data_log_force[ 926] <= 1'h0;
      write_done_data_log_force[ 927] <= 1'h0;
      write_done_data_log_force[ 928] <= 1'h0;
      write_done_data_log_force[ 929] <= 1'h0;
      write_done_data_log_force[ 930] <= 1'h0;
      write_done_data_log_force[ 931] <= 1'h0;
      write_done_data_log_force[ 932] <= 1'h0;
      write_done_data_log_force[ 933] <= 1'h0;
      write_done_data_log_force[ 934] <= 1'h0;
      write_done_data_log_force[ 935] <= 1'h0;
      write_done_data_log_force[ 936] <= 1'h0;
      write_done_data_log_force[ 937] <= 1'h0;
      write_done_data_log_force[ 938] <= 1'h0;
      write_done_data_log_force[ 939] <= 1'h0;
      write_done_data_log_force[ 940] <= 1'h0;
      write_done_data_log_force[ 941] <= 1'h0;
      write_done_data_log_force[ 942] <= 1'h0;
      write_done_data_log_force[ 943] <= 1'h0;
      write_done_data_log_force[ 944] <= 1'h0;
      write_done_data_log_force[ 945] <= 1'h0;
      write_done_data_log_force[ 946] <= 1'h0;
      write_done_data_log_force[ 947] <= 1'h0;
      write_done_data_log_force[ 948] <= 1'h0;
      write_done_data_log_force[ 949] <= 1'h0;
      write_done_data_log_force[ 950] <= 1'h0;
      write_done_data_log_force[ 951] <= 1'h0;
      write_done_data_log_force[ 952] <= 1'h0;
      write_done_data_log_force[ 953] <= 1'h0;
      write_done_data_log_force[ 954] <= 1'h0;
      write_done_data_log_force[ 955] <= 1'h0;
      write_done_data_log_force[ 956] <= 1'h0;
      write_done_data_log_force[ 957] <= 1'h0;
      write_done_data_log_force[ 958] <= 1'h0;
      write_done_data_log_force[ 959] <= 1'h0;
      write_done_data_log_force[ 960] <= 1'h0;
      write_done_data_log_force[ 961] <= 1'h0;
      write_done_data_log_force[ 962] <= 1'h0;
      write_done_data_log_force[ 963] <= 1'h0;
      write_done_data_log_force[ 964] <= 1'h0;
      write_done_data_log_force[ 965] <= 1'h0;
      write_done_data_log_force[ 966] <= 1'h0;
      write_done_data_log_force[ 967] <= 1'h0;
      write_done_data_log_force[ 968] <= 1'h0;
      write_done_data_log_force[ 969] <= 1'h0;
      write_done_data_log_force[ 970] <= 1'h0;
      write_done_data_log_force[ 971] <= 1'h0;
      write_done_data_log_force[ 972] <= 1'h0;
      write_done_data_log_force[ 973] <= 1'h0;
      write_done_data_log_force[ 974] <= 1'h0;
      write_done_data_log_force[ 975] <= 1'h0;
      write_done_data_log_force[ 976] <= 1'h0;
      write_done_data_log_force[ 977] <= 1'h0;
      write_done_data_log_force[ 978] <= 1'h0;
      write_done_data_log_force[ 979] <= 1'h0;
      write_done_data_log_force[ 980] <= 1'h0;
      write_done_data_log_force[ 981] <= 1'h0;
      write_done_data_log_force[ 982] <= 1'h0;
      write_done_data_log_force[ 983] <= 1'h0;
      write_done_data_log_force[ 984] <= 1'h0;
      write_done_data_log_force[ 985] <= 1'h0;
      write_done_data_log_force[ 986] <= 1'h0;
      write_done_data_log_force[ 987] <= 1'h0;
      write_done_data_log_force[ 988] <= 1'h0;
      write_done_data_log_force[ 989] <= 1'h0;
      write_done_data_log_force[ 990] <= 1'h0;
      write_done_data_log_force[ 991] <= 1'h0;
      write_done_data_log_force[ 992] <= 1'h0;
      write_done_data_log_force[ 993] <= 1'h0;
      write_done_data_log_force[ 994] <= 1'h0;
      write_done_data_log_force[ 995] <= 1'h0;
      write_done_data_log_force[ 996] <= 1'h0;
      write_done_data_log_force[ 997] <= 1'h0;
      write_done_data_log_force[ 998] <= 1'h0;
      write_done_data_log_force[ 999] <= 1'h0;
      write_done_data_log_force[1000] <= 1'h0;
      write_done_data_log_force[1001] <= 1'h0;
      write_done_data_log_force[1002] <= 1'h0;
      write_done_data_log_force[1003] <= 1'h0;
      write_done_data_log_force[1004] <= 1'h0;
      write_done_data_log_force[1005] <= 1'h0;
      write_done_data_log_force[1006] <= 1'h0;
      write_done_data_log_force[1007] <= 1'h0;
      write_done_data_log_force[1008] <= 1'h0;
      write_done_data_log_force[1009] <= 1'h0;
      write_done_data_log_force[1010] <= 1'h0;
      write_done_data_log_force[1011] <= 1'h0;
      write_done_data_log_force[1012] <= 1'h0;
      write_done_data_log_force[1013] <= 1'h0;
      write_done_data_log_force[1014] <= 1'h0;
      write_done_data_log_force[1015] <= 1'h0;
      write_done_data_log_force[1016] <= 1'h0;
      write_done_data_log_force[1017] <= 1'h0;
      write_done_data_log_force[1018] <= 1'h0;
      write_done_data_log_force[1019] <= 1'h0;
      write_done_data_log_force[1020] <= 1'h0;
      write_done_data_log_force[1021] <= 1'h0;
      write_done_data_log_force[1022] <= 1'h0;
      write_done_data_log_force[1023] <= 1'h0;
      write_done_data_log_force[1024] <= 1'h0;
      write_done_data_log_force[1025] <= 1'h0;
      write_done_data_log_force[1026] <= 1'h0;
      write_done_data_log_force[1027] <= 1'h0;
      write_done_data_log_force[1028] <= 1'h0;
      write_done_data_log_force[1029] <= 1'h0;
      write_done_data_log_force[1030] <= 1'h0;
      write_done_data_log_force[1031] <= 1'h0;
      write_done_data_log_force[1032] <= 1'h0;
      write_done_data_log_force[1033] <= 1'h0;
      write_done_data_log_force[1034] <= 1'h0;
      write_done_data_log_force[1035] <= 1'h0;
      write_done_data_log_force[1036] <= 1'h0;
      write_done_data_log_force[1037] <= 1'h0;
      write_done_data_log_force[1038] <= 1'h0;
      write_done_data_log_force[1039] <= 1'h0;
      write_done_data_log_force[1040] <= 1'h0;
      write_done_data_log_force[1041] <= 1'h0;
      write_done_data_log_force[1042] <= 1'h0;
      write_done_data_log_force[1043] <= 1'h0;
      write_done_data_log_force[1044] <= 1'h0;
      write_done_data_log_force[1045] <= 1'h0;
      write_done_data_log_force[1046] <= 1'h0;
      write_done_data_log_force[1047] <= 1'h0;
      write_done_data_log_force[1048] <= 1'h0;
      write_done_data_log_force[1049] <= 1'h0;
      write_done_data_log_force[1050] <= 1'h0;
      write_done_data_log_force[1051] <= 1'h0;
      write_done_data_log_force[1052] <= 1'h0;
      write_done_data_log_force[1053] <= 1'h0;
      write_done_data_log_force[1054] <= 1'h0;
      write_done_data_log_force[1055] <= 1'h0;
      write_done_data_log_force[1056] <= 1'h0;
      write_done_data_log_force[1057] <= 1'h0;
      write_done_data_log_force[1058] <= 1'h0;
      write_done_data_log_force[1059] <= 1'h0;
      write_done_data_log_force[1060] <= 1'h0;
      write_done_data_log_force[1061] <= 1'h0;
      write_done_data_log_force[1062] <= 1'h0;
      write_done_data_log_force[1063] <= 1'h0;
      write_done_data_log_force[1064] <= 1'h0;
      write_done_data_log_force[1065] <= 1'h0;
      write_done_data_log_force[1066] <= 1'h0;
      write_done_data_log_force[1067] <= 1'h0;
      write_done_data_log_force[1068] <= 1'h0;
      write_done_data_log_force[1069] <= 1'h0;
      write_done_data_log_force[1070] <= 1'h0;
      write_done_data_log_force[1071] <= 1'h0;
      write_done_data_log_force[1072] <= 1'h0;
      write_done_data_log_force[1073] <= 1'h0;
      write_done_data_log_force[1074] <= 1'h0;
      write_done_data_log_force[1075] <= 1'h0;
      write_done_data_log_force[1076] <= 1'h0;
      write_done_data_log_force[1077] <= 1'h0;
      write_done_data_log_force[1078] <= 1'h0;
      write_done_data_log_force[1079] <= 1'h0;
      write_done_data_log_force[1080] <= 1'h0;
      write_done_data_log_force[1081] <= 1'h0;
      write_done_data_log_force[1082] <= 1'h0;
      write_done_data_log_force[1083] <= 1'h0;
      write_done_data_log_force[1084] <= 1'h0;
      write_done_data_log_force[1085] <= 1'h0;
      write_done_data_log_force[1086] <= 1'h0;
      write_done_data_log_force[1087] <= 1'h0;
      write_done_data_log_force[1088] <= 1'h0;
      write_done_data_log_force[1089] <= 1'h0;
      write_done_data_log_force[1090] <= 1'h0;
      write_done_data_log_force[1091] <= 1'h0;
      write_done_data_log_force[1092] <= 1'h0;
      write_done_data_log_force[1093] <= 1'h0;
      write_done_data_log_force[1094] <= 1'h0;
      write_done_data_log_force[1095] <= 1'h0;
      write_done_data_log_force[1096] <= 1'h0;
      write_done_data_log_force[1097] <= 1'h0;
      write_done_data_log_force[1098] <= 1'h0;
      write_done_data_log_force[1099] <= 1'h0;
      write_done_data_log_force[1100] <= 1'h0;
      write_done_data_log_force[1101] <= 1'h0;
      write_done_data_log_force[1102] <= 1'h0;
      write_done_data_log_force[1103] <= 1'h0;
      write_done_data_log_force[1104] <= 1'h0;
      write_done_data_log_force[1105] <= 1'h0;
      write_done_data_log_force[1106] <= 1'h0;
      write_done_data_log_force[1107] <= 1'h0;
      write_done_data_log_force[1108] <= 1'h0;
      write_done_data_log_force[1109] <= 1'h0;
      write_done_data_log_force[1110] <= 1'h0;
      write_done_data_log_force[1111] <= 1'h0;
      write_done_data_log_force[1112] <= 1'h0;
      write_done_data_log_force[1113] <= 1'h0;
      write_done_data_log_force[1114] <= 1'h0;
      write_done_data_log_force[1115] <= 1'h0;
      write_done_data_log_force[1116] <= 1'h0;
      write_done_data_log_force[1117] <= 1'h0;
      write_done_data_log_force[1118] <= 1'h0;
      write_done_data_log_force[1119] <= 1'h0;
      write_done_data_log_force[1120] <= 1'h0;
      write_done_data_log_force[1121] <= 1'h0;
      write_done_data_log_force[1122] <= 1'h0;
      write_done_data_log_force[1123] <= 1'h0;
      write_done_data_log_force[1124] <= 1'h0;
      write_done_data_log_force[1125] <= 1'h0;
      write_done_data_log_force[1126] <= 1'h0;
      write_done_data_log_force[1127] <= 1'h0;
      write_done_data_log_force[1128] <= 1'h0;
      write_done_data_log_force[1129] <= 1'h0;
      write_done_data_log_force[1130] <= 1'h0;
      write_done_data_log_force[1131] <= 1'h0;
      write_done_data_log_force[1132] <= 1'h0;
      write_done_data_log_force[1133] <= 1'h0;
      write_done_data_log_force[1134] <= 1'h0;
      write_done_data_log_force[1135] <= 1'h0;
      write_done_data_log_force[1136] <= 1'h0;
      write_done_data_log_force[1137] <= 1'h0;
      write_done_data_log_force[1138] <= 1'h0;
      write_done_data_log_force[1139] <= 1'h0;
      write_done_data_log_force[1140] <= 1'h0;
      write_done_data_log_force[1141] <= 1'h0;
      write_done_data_log_force[1142] <= 1'h0;
      write_done_data_log_force[1143] <= 1'h0;
      write_done_data_log_force[1144] <= 1'h0;
      write_done_data_log_force[1145] <= 1'h0;
      write_done_data_log_force[1146] <= 1'h0;
      write_done_data_log_force[1147] <= 1'h0;
      write_done_data_log_force[1148] <= 1'h0;
      write_done_data_log_force[1149] <= 1'h0;
      write_done_data_log_force[1150] <= 1'h0;
      write_done_data_log_force[1151] <= 1'h0;
      write_done_data_log_force[1152] <= 1'h0;
      write_done_data_log_force[1153] <= 1'h0;
      write_done_data_log_force[1154] <= 1'h0;
      write_done_data_log_force[1155] <= 1'h0;
      write_done_data_log_force[1156] <= 1'h0;
      write_done_data_log_force[1157] <= 1'h0;
      write_done_data_log_force[1158] <= 1'h0;
      write_done_data_log_force[1159] <= 1'h0;
      write_done_data_log_force[1160] <= 1'h0;
      write_done_data_log_force[1161] <= 1'h0;
      write_done_data_log_force[1162] <= 1'h0;
      write_done_data_log_force[1163] <= 1'h0;
      write_done_data_log_force[1164] <= 1'h0;
      write_done_data_log_force[1165] <= 1'h0;
      write_done_data_log_force[1166] <= 1'h0;
      write_done_data_log_force[1167] <= 1'h0;
      write_done_data_log_force[1168] <= 1'h0;
      write_done_data_log_force[1169] <= 1'h0;
      write_done_data_log_force[1170] <= 1'h0;
      write_done_data_log_force[1171] <= 1'h0;
      write_done_data_log_force[1172] <= 1'h0;
      write_done_data_log_force[1173] <= 1'h0;
      write_done_data_log_force[1174] <= 1'h0;
      write_done_data_log_force[1175] <= 1'h0;
      write_done_data_log_force[1176] <= 1'h0;
      write_done_data_log_force[1177] <= 1'h0;
      write_done_data_log_force[1178] <= 1'h0;
      write_done_data_log_force[1179] <= 1'h0;
      write_done_data_log_force[1180] <= 1'h0;
      write_done_data_log_force[1181] <= 1'h0;
      write_done_data_log_force[1182] <= 1'h0;
      write_done_data_log_force[1183] <= 1'h0;
      write_done_data_log_force[1184] <= 1'h0;
      write_done_data_log_force[1185] <= 1'h0;
      write_done_data_log_force[1186] <= 1'h0;
      write_done_data_log_force[1187] <= 1'h0;
      write_done_data_log_force[1188] <= 1'h0;
      write_done_data_log_force[1189] <= 1'h0;
      write_done_data_log_force[1190] <= 1'h0;
      write_done_data_log_force[1191] <= 1'h0;
      write_done_data_log_force[1192] <= 1'h0;
      write_done_data_log_force[1193] <= 1'h0;
      write_done_data_log_force[1194] <= 1'h0;
      write_done_data_log_force[1195] <= 1'h0;
      write_done_data_log_force[1196] <= 1'h0;
      write_done_data_log_force[1197] <= 1'h0;
      write_done_data_log_force[1198] <= 1'h0;
      write_done_data_log_force[1199] <= 1'h0;
      write_done_data_log_force[1200] <= 1'h0;
      write_done_data_log_force[1201] <= 1'h0;
      write_done_data_log_force[1202] <= 1'h0;
      write_done_data_log_force[1203] <= 1'h0;
      write_done_data_log_force[1204] <= 1'h0;
      write_done_data_log_force[1205] <= 1'h0;
      write_done_data_log_force[1206] <= 1'h0;
      write_done_data_log_force[1207] <= 1'h0;
      write_done_data_log_force[1208] <= 1'h0;
      write_done_data_log_force[1209] <= 1'h0;
      write_done_data_log_force[1210] <= 1'h0;
      write_done_data_log_force[1211] <= 1'h0;
      write_done_data_log_force[1212] <= 1'h0;
      write_done_data_log_force[1213] <= 1'h0;
      write_done_data_log_force[1214] <= 1'h0;
      write_done_data_log_force[1215] <= 1'h0;
      write_done_data_log_force[1216] <= 1'h0;
      write_done_data_log_force[1217] <= 1'h0;
      write_done_data_log_force[1218] <= 1'h0;
      write_done_data_log_force[1219] <= 1'h0;
      write_done_data_log_force[1220] <= 1'h0;
      write_done_data_log_force[1221] <= 1'h0;
      write_done_data_log_force[1222] <= 1'h0;
      write_done_data_log_force[1223] <= 1'h0;
      write_done_data_log_force[1224] <= 1'h0;
      write_done_data_log_force[1225] <= 1'h0;
      write_done_data_log_force[1226] <= 1'h0;
      write_done_data_log_force[1227] <= 1'h0;
      write_done_data_log_force[1228] <= 1'h0;
      write_done_data_log_force[1229] <= 1'h0;
      write_done_data_log_force[1230] <= 1'h0;
      write_done_data_log_force[1231] <= 1'h0;
      write_done_data_log_force[1232] <= 1'h0;
      write_done_data_log_force[1233] <= 1'h0;
      write_done_data_log_force[1234] <= 1'h0;
      write_done_data_log_force[1235] <= 1'h0;
      write_done_data_log_force[1236] <= 1'h0;
      write_done_data_log_force[1237] <= 1'h0;
      write_done_data_log_force[1238] <= 1'h0;
      write_done_data_log_force[1239] <= 1'h0;
      write_done_data_log_force[1240] <= 1'h0;
      write_done_data_log_force[1241] <= 1'h0;
      write_done_data_log_force[1242] <= 1'h0;
      write_done_data_log_force[1243] <= 1'h0;
      write_done_data_log_force[1244] <= 1'h0;
      write_done_data_log_force[1245] <= 1'h0;
      write_done_data_log_force[1246] <= 1'h0;
      write_done_data_log_force[1247] <= 1'h0;
      write_done_data_log_force[1248] <= 1'h0;
      write_done_data_log_force[1249] <= 1'h0;
      write_done_data_log_force[1250] <= 1'h0;
      write_done_data_log_force[1251] <= 1'h0;
      write_done_data_log_force[1252] <= 1'h0;
      write_done_data_log_force[1253] <= 1'h0;
      write_done_data_log_force[1254] <= 1'h0;
      write_done_data_log_force[1255] <= 1'h0;
      write_done_data_log_force[1256] <= 1'h0;
      write_done_data_log_force[1257] <= 1'h0;
      write_done_data_log_force[1258] <= 1'h0;
      write_done_data_log_force[1259] <= 1'h0;
      write_done_data_log_force[1260] <= 1'h0;
      write_done_data_log_force[1261] <= 1'h0;
      write_done_data_log_force[1262] <= 1'h0;
      write_done_data_log_force[1263] <= 1'h0;
      write_done_data_log_force[1264] <= 1'h0;
      write_done_data_log_force[1265] <= 1'h0;
      write_done_data_log_force[1266] <= 1'h0;
      write_done_data_log_force[1267] <= 1'h0;
      write_done_data_log_force[1268] <= 1'h0;
      write_done_data_log_force[1269] <= 1'h0;
      write_done_data_log_force[1270] <= 1'h0;
      write_done_data_log_force[1271] <= 1'h0;
      write_done_data_log_force[1272] <= 1'h0;
      write_done_data_log_force[1273] <= 1'h0;
      write_done_data_log_force[1274] <= 1'h0;
      write_done_data_log_force[1275] <= 1'h0;
      write_done_data_log_force[1276] <= 1'h0;
      write_done_data_log_force[1277] <= 1'h0;
      write_done_data_log_force[1278] <= 1'h0;
      write_done_data_log_force[1279] <= 1'h0;
      write_done_data_log_force[1280] <= 1'h0;
      write_done_data_log_force[1281] <= 1'h0;
      write_done_data_log_force[1282] <= 1'h0;
      write_done_data_log_force[1283] <= 1'h0;
      write_done_data_log_force[1284] <= 1'h0;
      write_done_data_log_force[1285] <= 1'h0;
      write_done_data_log_force[1286] <= 1'h0;
      write_done_data_log_force[1287] <= 1'h0;
      write_done_data_log_force[1288] <= 1'h0;
      write_done_data_log_force[1289] <= 1'h0;
      write_done_data_log_force[1290] <= 1'h0;
      write_done_data_log_force[1291] <= 1'h0;
      write_done_data_log_force[1292] <= 1'h0;
      write_done_data_log_force[1293] <= 1'h0;
      write_done_data_log_force[1294] <= 1'h0;
      write_done_data_log_force[1295] <= 1'h0;
      write_done_data_log_force[1296] <= 1'h0;
      write_done_data_log_force[1297] <= 1'h0;
      write_done_data_log_force[1298] <= 1'h0;
      write_done_data_log_force[1299] <= 1'h0;
      write_done_data_log_force[1300] <= 1'h0;
      write_done_data_log_force[1301] <= 1'h0;
      write_done_data_log_force[1302] <= 1'h0;
      write_done_data_log_force[1303] <= 1'h0;
      write_done_data_log_force[1304] <= 1'h0;
      write_done_data_log_force[1305] <= 1'h0;
      write_done_data_log_force[1306] <= 1'h0;
      write_done_data_log_force[1307] <= 1'h0;
      write_done_data_log_force[1308] <= 1'h0;
      write_done_data_log_force[1309] <= 1'h0;
      write_done_data_log_force[1310] <= 1'h0;
      write_done_data_log_force[1311] <= 1'h0;
      write_done_data_log_force[1312] <= 1'h0;
      write_done_data_log_force[1313] <= 1'h0;
      write_done_data_log_force[1314] <= 1'h0;
      write_done_data_log_force[1315] <= 1'h0;
      write_done_data_log_force[1316] <= 1'h0;
      write_done_data_log_force[1317] <= 1'h0;
      write_done_data_log_force[1318] <= 1'h0;
      write_done_data_log_force[1319] <= 1'h0;
      write_done_data_log_force[1320] <= 1'h0;
      write_done_data_log_force[1321] <= 1'h0;
      write_done_data_log_force[1322] <= 1'h0;
      write_done_data_log_force[1323] <= 1'h0;
      write_done_data_log_force[1324] <= 1'h0;
      write_done_data_log_force[1325] <= 1'h0;
      write_done_data_log_force[1326] <= 1'h0;
      write_done_data_log_force[1327] <= 1'h0;
      write_done_data_log_force[1328] <= 1'h0;
      write_done_data_log_force[1329] <= 1'h0;
      write_done_data_log_force[1330] <= 1'h0;
      write_done_data_log_force[1331] <= 1'h0;
      write_done_data_log_force[1332] <= 1'h0;
      write_done_data_log_force[1333] <= 1'h0;
      write_done_data_log_force[1334] <= 1'h0;
      write_done_data_log_force[1335] <= 1'h0;
      write_done_data_log_force[1336] <= 1'h0;
      write_done_data_log_force[1337] <= 1'h0;
      write_done_data_log_force[1338] <= 1'h0;
      write_done_data_log_force[1339] <= 1'h0;
      write_done_data_log_force[1340] <= 1'h0;
      write_done_data_log_force[1341] <= 1'h0;
      write_done_data_log_force[1342] <= 1'h0;
      write_done_data_log_force[1343] <= 1'h0;
      write_done_data_log_force[1344] <= 1'h0;
      write_done_data_log_force[1345] <= 1'h0;
      write_done_data_log_force[1346] <= 1'h0;
      write_done_data_log_force[1347] <= 1'h0;
      write_done_data_log_force[1348] <= 1'h0;
      write_done_data_log_force[1349] <= 1'h0;
      write_done_data_log_force[1350] <= 1'h0;
      write_done_data_log_force[1351] <= 1'h0;
      write_done_data_log_force[1352] <= 1'h0;
      write_done_data_log_force[1353] <= 1'h0;
      write_done_data_log_force[1354] <= 1'h0;
      write_done_data_log_force[1355] <= 1'h0;
      write_done_data_log_force[1356] <= 1'h0;
      write_done_data_log_force[1357] <= 1'h0;
      write_done_data_log_force[1358] <= 1'h0;
      write_done_data_log_force[1359] <= 1'h0;
      write_done_data_log_force[1360] <= 1'h0;
      write_done_data_log_force[1361] <= 1'h0;
      write_done_data_log_force[1362] <= 1'h0;
      write_done_data_log_force[1363] <= 1'h0;
      write_done_data_log_force[1364] <= 1'h0;
      write_done_data_log_force[1365] <= 1'h0;
      write_done_data_log_force[1366] <= 1'h0;
      write_done_data_log_force[1367] <= 1'h0;
      write_done_data_log_force[1368] <= 1'h0;
      write_done_data_log_force[1369] <= 1'h0;
      write_done_data_log_force[1370] <= 1'h0;
      write_done_data_log_force[1371] <= 1'h0;
      write_done_data_log_force[1372] <= 1'h0;
      write_done_data_log_force[1373] <= 1'h0;
      write_done_data_log_force[1374] <= 1'h0;
      write_done_data_log_force[1375] <= 1'h0;
      write_done_data_log_force[1376] <= 1'h0;
      write_done_data_log_force[1377] <= 1'h0;
      write_done_data_log_force[1378] <= 1'h0;
      write_done_data_log_force[1379] <= 1'h0;
      write_done_data_log_force[1380] <= 1'h0;
      write_done_data_log_force[1381] <= 1'h0;
      write_done_data_log_force[1382] <= 1'h0;
      write_done_data_log_force[1383] <= 1'h0;
      write_done_data_log_force[1384] <= 1'h0;
      write_done_data_log_force[1385] <= 1'h0;
      write_done_data_log_force[1386] <= 1'h0;
      write_done_data_log_force[1387] <= 1'h0;
      write_done_data_log_force[1388] <= 1'h0;
      write_done_data_log_force[1389] <= 1'h0;
      write_done_data_log_force[1390] <= 1'h0;
      write_done_data_log_force[1391] <= 1'h0;
      write_done_data_log_force[1392] <= 1'h0;
      write_done_data_log_force[1393] <= 1'h0;
      write_done_data_log_force[1394] <= 1'h0;
      write_done_data_log_force[1395] <= 1'h0;
      write_done_data_log_force[1396] <= 1'h0;
      write_done_data_log_force[1397] <= 1'h0;
      write_done_data_log_force[1398] <= 1'h0;
      write_done_data_log_force[1399] <= 1'h0;
      write_done_data_log_force[1400] <= 1'h0;
      write_done_data_log_force[1401] <= 1'h0;
      write_done_data_log_force[1402] <= 1'h0;
      write_done_data_log_force[1403] <= 1'h0;
      write_done_data_log_force[1404] <= 1'h0;
      write_done_data_log_force[1405] <= 1'h0;
      write_done_data_log_force[1406] <= 1'h0;
      write_done_data_log_force[1407] <= 1'h0;
      write_done_data_log_force[1408] <= 1'h0;
      write_done_data_log_force[1409] <= 1'h0;
      write_done_data_log_force[1410] <= 1'h0;
      write_done_data_log_force[1411] <= 1'h0;
      write_done_data_log_force[1412] <= 1'h0;
      write_done_data_log_force[1413] <= 1'h0;
      write_done_data_log_force[1414] <= 1'h0;
      write_done_data_log_force[1415] <= 1'h0;
      write_done_data_log_force[1416] <= 1'h0;
      write_done_data_log_force[1417] <= 1'h0;
      write_done_data_log_force[1418] <= 1'h0;
      write_done_data_log_force[1419] <= 1'h0;
      write_done_data_log_force[1420] <= 1'h0;
      write_done_data_log_force[1421] <= 1'h0;
      write_done_data_log_force[1422] <= 1'h0;
      write_done_data_log_force[1423] <= 1'h0;
      write_done_data_log_force[1424] <= 1'h0;
      write_done_data_log_force[1425] <= 1'h0;
      write_done_data_log_force[1426] <= 1'h0;
      write_done_data_log_force[1427] <= 1'h0;
      write_done_data_log_force[1428] <= 1'h0;
      write_done_data_log_force[1429] <= 1'h0;
      write_done_data_log_force[1430] <= 1'h0;
      write_done_data_log_force[1431] <= 1'h0;
      write_done_data_log_force[1432] <= 1'h0;
      write_done_data_log_force[1433] <= 1'h0;
      write_done_data_log_force[1434] <= 1'h0;
      write_done_data_log_force[1435] <= 1'h0;
      write_done_data_log_force[1436] <= 1'h0;
      write_done_data_log_force[1437] <= 1'h0;
      write_done_data_log_force[1438] <= 1'h0;
      write_done_data_log_force[1439] <= 1'h0;
      write_done_data_log_force[1440] <= 1'h0;
      write_done_data_log_force[1441] <= 1'h0;
      write_done_data_log_force[1442] <= 1'h0;
      write_done_data_log_force[1443] <= 1'h0;
      write_done_data_log_force[1444] <= 1'h0;
      write_done_data_log_force[1445] <= 1'h0;
      write_done_data_log_force[1446] <= 1'h0;
      write_done_data_log_force[1447] <= 1'h0;
      write_done_data_log_force[1448] <= 1'h0;
      write_done_data_log_force[1449] <= 1'h0;
      write_done_data_log_force[1450] <= 1'h0;
      write_done_data_log_force[1451] <= 1'h0;
      write_done_data_log_force[1452] <= 1'h0;
      write_done_data_log_force[1453] <= 1'h0;
      write_done_data_log_force[1454] <= 1'h0;
      write_done_data_log_force[1455] <= 1'h0;
      write_done_data_log_force[1456] <= 1'h0;
      write_done_data_log_force[1457] <= 1'h0;
      write_done_data_log_force[1458] <= 1'h0;
      write_done_data_log_force[1459] <= 1'h0;
      write_done_data_log_force[1460] <= 1'h0;
      write_done_data_log_force[1461] <= 1'h0;
      write_done_data_log_force[1462] <= 1'h0;
      write_done_data_log_force[1463] <= 1'h0;
      write_done_data_log_force[1464] <= 1'h0;
      write_done_data_log_force[1465] <= 1'h0;
      write_done_data_log_force[1466] <= 1'h0;
      write_done_data_log_force[1467] <= 1'h0;
      write_done_data_log_force[1468] <= 1'h0;
      write_done_data_log_force[1469] <= 1'h0;
      write_done_data_log_force[1470] <= 1'h0;
      write_done_data_log_force[1471] <= 1'h0;
      write_done_data_log_force[1472] <= 1'h0;
      write_done_data_log_force[1473] <= 1'h0;
      write_done_data_log_force[1474] <= 1'h0;
      write_done_data_log_force[1475] <= 1'h0;
      write_done_data_log_force[1476] <= 1'h0;
      write_done_data_log_force[1477] <= 1'h0;
      write_done_data_log_force[1478] <= 1'h0;
      write_done_data_log_force[1479] <= 1'h0;
      write_done_data_log_force[1480] <= 1'h0;
      write_done_data_log_force[1481] <= 1'h0;
      write_done_data_log_force[1482] <= 1'h0;
      write_done_data_log_force[1483] <= 1'h0;
      write_done_data_log_force[1484] <= 1'h0;
      write_done_data_log_force[1485] <= 1'h0;
      write_done_data_log_force[1486] <= 1'h0;
      write_done_data_log_force[1487] <= 1'h0;
      write_done_data_log_force[1488] <= 1'h0;
      write_done_data_log_force[1489] <= 1'h0;
      write_done_data_log_force[1490] <= 1'h0;
      write_done_data_log_force[1491] <= 1'h0;
      write_done_data_log_force[1492] <= 1'h0;
      write_done_data_log_force[1493] <= 1'h0;
      write_done_data_log_force[1494] <= 1'h0;
      write_done_data_log_force[1495] <= 1'h0;
      write_done_data_log_force[1496] <= 1'h0;
      write_done_data_log_force[1497] <= 1'h0;
      write_done_data_log_force[1498] <= 1'h0;
      write_done_data_log_force[1499] <= 1'h0;
      write_done_data_log_force[1500] <= 1'h0;
      write_done_data_log_force[1501] <= 1'h0;
      write_done_data_log_force[1502] <= 1'h0;
      write_done_data_log_force[1503] <= 1'h0;
      write_done_data_log_force[1504] <= 1'h0;
      write_done_data_log_force[1505] <= 1'h0;
      write_done_data_log_force[1506] <= 1'h0;
      write_done_data_log_force[1507] <= 1'h0;
      write_done_data_log_force[1508] <= 1'h0;
      write_done_data_log_force[1509] <= 1'h0;
      write_done_data_log_force[1510] <= 1'h0;
      write_done_data_log_force[1511] <= 1'h0;
      write_done_data_log_force[1512] <= 1'h0;
      write_done_data_log_force[1513] <= 1'h0;
      write_done_data_log_force[1514] <= 1'h0;
      write_done_data_log_force[1515] <= 1'h0;
      write_done_data_log_force[1516] <= 1'h0;
      write_done_data_log_force[1517] <= 1'h0;
      write_done_data_log_force[1518] <= 1'h0;
      write_done_data_log_force[1519] <= 1'h0;
      write_done_data_log_force[1520] <= 1'h0;
      write_done_data_log_force[1521] <= 1'h0;
      write_done_data_log_force[1522] <= 1'h0;
      write_done_data_log_force[1523] <= 1'h0;
      write_done_data_log_force[1524] <= 1'h0;
      write_done_data_log_force[1525] <= 1'h0;
      write_done_data_log_force[1526] <= 1'h0;
      write_done_data_log_force[1527] <= 1'h0;
      write_done_data_log_force[1528] <= 1'h0;
      write_done_data_log_force[1529] <= 1'h0;
      write_done_data_log_force[1530] <= 1'h0;
      write_done_data_log_force[1531] <= 1'h0;
      write_done_data_log_force[1532] <= 1'h0;
      write_done_data_log_force[1533] <= 1'h0;
      write_done_data_log_force[1534] <= 1'h0;
      write_done_data_log_force[1535] <= 1'h0;
      write_done_data_log_force[1536] <= 1'h0;
      write_done_data_log_force[1537] <= 1'h0;
      write_done_data_log_force[1538] <= 1'h0;
      write_done_data_log_force[1539] <= 1'h0;
      write_done_data_log_force[1540] <= 1'h0;
      write_done_data_log_force[1541] <= 1'h0;
      write_done_data_log_force[1542] <= 1'h0;
      write_done_data_log_force[1543] <= 1'h0;
      write_done_data_log_force[1544] <= 1'h0;
      write_done_data_log_force[1545] <= 1'h0;
      write_done_data_log_force[1546] <= 1'h0;
      write_done_data_log_force[1547] <= 1'h0;
      write_done_data_log_force[1548] <= 1'h0;
      write_done_data_log_force[1549] <= 1'h0;
      write_done_data_log_force[1550] <= 1'h0;
      write_done_data_log_force[1551] <= 1'h0;
      write_done_data_log_force[1552] <= 1'h0;
      write_done_data_log_force[1553] <= 1'h0;
      write_done_data_log_force[1554] <= 1'h0;
      write_done_data_log_force[1555] <= 1'h0;
      write_done_data_log_force[1556] <= 1'h0;
      write_done_data_log_force[1557] <= 1'h0;
      write_done_data_log_force[1558] <= 1'h0;
      write_done_data_log_force[1559] <= 1'h0;
      write_done_data_log_force[1560] <= 1'h0;
      write_done_data_log_force[1561] <= 1'h0;
      write_done_data_log_force[1562] <= 1'h0;
      write_done_data_log_force[1563] <= 1'h0;
      write_done_data_log_force[1564] <= 1'h0;
      write_done_data_log_force[1565] <= 1'h0;
      write_done_data_log_force[1566] <= 1'h0;
      write_done_data_log_force[1567] <= 1'h0;
      write_done_data_log_force[1568] <= 1'h0;
      write_done_data_log_force[1569] <= 1'h0;
      write_done_data_log_force[1570] <= 1'h0;
      write_done_data_log_force[1571] <= 1'h0;
      write_done_data_log_force[1572] <= 1'h0;
      write_done_data_log_force[1573] <= 1'h0;
      write_done_data_log_force[1574] <= 1'h0;
      write_done_data_log_force[1575] <= 1'h0;
      write_done_data_log_force[1576] <= 1'h0;
      write_done_data_log_force[1577] <= 1'h0;
      write_done_data_log_force[1578] <= 1'h0;
      write_done_data_log_force[1579] <= 1'h0;
      write_done_data_log_force[1580] <= 1'h0;
      write_done_data_log_force[1581] <= 1'h0;
      write_done_data_log_force[1582] <= 1'h0;
      write_done_data_log_force[1583] <= 1'h0;
      write_done_data_log_force[1584] <= 1'h0;
      write_done_data_log_force[1585] <= 1'h0;
      write_done_data_log_force[1586] <= 1'h0;
      write_done_data_log_force[1587] <= 1'h0;
      write_done_data_log_force[1588] <= 1'h0;
      write_done_data_log_force[1589] <= 1'h0;
      write_done_data_log_force[1590] <= 1'h0;
      write_done_data_log_force[1591] <= 1'h0;
      write_done_data_log_force[1592] <= 1'h0;
      write_done_data_log_force[1593] <= 1'h0;
      write_done_data_log_force[1594] <= 1'h0;
      write_done_data_log_force[1595] <= 1'h0;
      write_done_data_log_force[1596] <= 1'h0;
      write_done_data_log_force[1597] <= 1'h0;
      write_done_data_log_force[1598] <= 1'h0;
      write_done_data_log_force[1599] <= 1'h0;
      write_done_data_log_force[1600] <= 1'h0;
      write_done_data_log_force[1601] <= 1'h0;
      write_done_data_log_force[1602] <= 1'h0;
      write_done_data_log_force[1603] <= 1'h0;
      write_done_data_log_force[1604] <= 1'h0;
      write_done_data_log_force[1605] <= 1'h0;
      write_done_data_log_force[1606] <= 1'h0;
      write_done_data_log_force[1607] <= 1'h0;
      write_done_data_log_force[1608] <= 1'h0;
      write_done_data_log_force[1609] <= 1'h0;
      write_done_data_log_force[1610] <= 1'h0;
      write_done_data_log_force[1611] <= 1'h0;
      write_done_data_log_force[1612] <= 1'h0;
      write_done_data_log_force[1613] <= 1'h0;
      write_done_data_log_force[1614] <= 1'h0;
      write_done_data_log_force[1615] <= 1'h0;
      write_done_data_log_force[1616] <= 1'h0;
      write_done_data_log_force[1617] <= 1'h0;
      write_done_data_log_force[1618] <= 1'h0;
      write_done_data_log_force[1619] <= 1'h0;
      write_done_data_log_force[1620] <= 1'h0;
      write_done_data_log_force[1621] <= 1'h0;
      write_done_data_log_force[1622] <= 1'h0;
      write_done_data_log_force[1623] <= 1'h0;
      write_done_data_log_force[1624] <= 1'h0;
      write_done_data_log_force[1625] <= 1'h0;
      write_done_data_log_force[1626] <= 1'h0;
      write_done_data_log_force[1627] <= 1'h0;
      write_done_data_log_force[1628] <= 1'h0;
      write_done_data_log_force[1629] <= 1'h0;
      write_done_data_log_force[1630] <= 1'h0;
      write_done_data_log_force[1631] <= 1'h0;
      write_done_data_log_force[1632] <= 1'h0;
      write_done_data_log_force[1633] <= 1'h0;
      write_done_data_log_force[1634] <= 1'h0;
      write_done_data_log_force[1635] <= 1'h0;
      write_done_data_log_force[1636] <= 1'h0;
      write_done_data_log_force[1637] <= 1'h0;
      write_done_data_log_force[1638] <= 1'h0;
      write_done_data_log_force[1639] <= 1'h0;
      write_done_data_log_force[1640] <= 1'h0;
      write_done_data_log_force[1641] <= 1'h0;
      write_done_data_log_force[1642] <= 1'h0;
      write_done_data_log_force[1643] <= 1'h0;
      write_done_data_log_force[1644] <= 1'h0;
      write_done_data_log_force[1645] <= 1'h0;
      write_done_data_log_force[1646] <= 1'h0;
      write_done_data_log_force[1647] <= 1'h0;
      write_done_data_log_force[1648] <= 1'h0;
      write_done_data_log_force[1649] <= 1'h0;
      write_done_data_log_force[1650] <= 1'h0;
      write_done_data_log_force[1651] <= 1'h0;
      write_done_data_log_force[1652] <= 1'h0;
      write_done_data_log_force[1653] <= 1'h0;
      write_done_data_log_force[1654] <= 1'h0;
      write_done_data_log_force[1655] <= 1'h0;
      write_done_data_log_force[1656] <= 1'h0;
      write_done_data_log_force[1657] <= 1'h0;
      write_done_data_log_force[1658] <= 1'h0;
      write_done_data_log_force[1659] <= 1'h0;
      write_done_data_log_force[1660] <= 1'h0;
      write_done_data_log_force[1661] <= 1'h0;
      write_done_data_log_force[1662] <= 1'h0;
      write_done_data_log_force[1663] <= 1'h0;
      write_done_data_log_force[1664] <= 1'h0;
      write_done_data_log_force[1665] <= 1'h0;
      write_done_data_log_force[1666] <= 1'h0;
      write_done_data_log_force[1667] <= 1'h0;
      write_done_data_log_force[1668] <= 1'h0;
      write_done_data_log_force[1669] <= 1'h0;
      write_done_data_log_force[1670] <= 1'h0;
      write_done_data_log_force[1671] <= 1'h0;
      write_done_data_log_force[1672] <= 1'h0;
      write_done_data_log_force[1673] <= 1'h0;
      write_done_data_log_force[1674] <= 1'h0;
      write_done_data_log_force[1675] <= 1'h0;
      write_done_data_log_force[1676] <= 1'h0;
      write_done_data_log_force[1677] <= 1'h0;
      write_done_data_log_force[1678] <= 1'h0;
      write_done_data_log_force[1679] <= 1'h0;
      write_done_data_log_force[1680] <= 1'h0;
      write_done_data_log_force[1681] <= 1'h0;
      write_done_data_log_force[1682] <= 1'h0;
      write_done_data_log_force[1683] <= 1'h0;
      write_done_data_log_force[1684] <= 1'h0;
      write_done_data_log_force[1685] <= 1'h0;
      write_done_data_log_force[1686] <= 1'h0;
      write_done_data_log_force[1687] <= 1'h0;
      write_done_data_log_force[1688] <= 1'h0;
      write_done_data_log_force[1689] <= 1'h0;
      write_done_data_log_force[1690] <= 1'h0;
      write_done_data_log_force[1691] <= 1'h0;
      write_done_data_log_force[1692] <= 1'h0;
      write_done_data_log_force[1693] <= 1'h0;
      write_done_data_log_force[1694] <= 1'h0;
      write_done_data_log_force[1695] <= 1'h0;
      write_done_data_log_force[1696] <= 1'h0;
      write_done_data_log_force[1697] <= 1'h0;
      write_done_data_log_force[1698] <= 1'h0;
      write_done_data_log_force[1699] <= 1'h0;
      write_done_data_log_force[1700] <= 1'h0;
      write_done_data_log_force[1701] <= 1'h0;
      write_done_data_log_force[1702] <= 1'h0;
      write_done_data_log_force[1703] <= 1'h0;
      write_done_data_log_force[1704] <= 1'h0;
      write_done_data_log_force[1705] <= 1'h0;
      write_done_data_log_force[1706] <= 1'h0;
      write_done_data_log_force[1707] <= 1'h0;
      write_done_data_log_force[1708] <= 1'h0;
      write_done_data_log_force[1709] <= 1'h0;
      write_done_data_log_force[1710] <= 1'h0;
      write_done_data_log_force[1711] <= 1'h0;
      write_done_data_log_force[1712] <= 1'h0;
      write_done_data_log_force[1713] <= 1'h0;
      write_done_data_log_force[1714] <= 1'h0;
      write_done_data_log_force[1715] <= 1'h0;
      write_done_data_log_force[1716] <= 1'h0;
      write_done_data_log_force[1717] <= 1'h0;
      write_done_data_log_force[1718] <= 1'h0;
      write_done_data_log_force[1719] <= 1'h0;
      write_done_data_log_force[1720] <= 1'h0;
      write_done_data_log_force[1721] <= 1'h0;
      write_done_data_log_force[1722] <= 1'h0;
      write_done_data_log_force[1723] <= 1'h0;
      write_done_data_log_force[1724] <= 1'h0;
      write_done_data_log_force[1725] <= 1'h0;
      write_done_data_log_force[1726] <= 1'h0;
      write_done_data_log_force[1727] <= 1'h0;
      write_done_data_log_force[1728] <= 1'h0;
      write_done_data_log_force[1729] <= 1'h0;
      write_done_data_log_force[1730] <= 1'h0;
      write_done_data_log_force[1731] <= 1'h0;
      write_done_data_log_force[1732] <= 1'h0;
      write_done_data_log_force[1733] <= 1'h0;
      write_done_data_log_force[1734] <= 1'h0;
      write_done_data_log_force[1735] <= 1'h0;
      write_done_data_log_force[1736] <= 1'h0;
      write_done_data_log_force[1737] <= 1'h0;
      write_done_data_log_force[1738] <= 1'h0;
      write_done_data_log_force[1739] <= 1'h0;
      write_done_data_log_force[1740] <= 1'h0;
      write_done_data_log_force[1741] <= 1'h0;
      write_done_data_log_force[1742] <= 1'h0;
      write_done_data_log_force[1743] <= 1'h0;
      write_done_data_log_force[1744] <= 1'h0;
      write_done_data_log_force[1745] <= 1'h0;
      write_done_data_log_force[1746] <= 1'h0;
      write_done_data_log_force[1747] <= 1'h0;
      write_done_data_log_force[1748] <= 1'h0;
      write_done_data_log_force[1749] <= 1'h0;
      write_done_data_log_force[1750] <= 1'h0;
      write_done_data_log_force[1751] <= 1'h0;
      write_done_data_log_force[1752] <= 1'h0;
      write_done_data_log_force[1753] <= 1'h0;
      write_done_data_log_force[1754] <= 1'h0;
      write_done_data_log_force[1755] <= 1'h0;
      write_done_data_log_force[1756] <= 1'h0;
      write_done_data_log_force[1757] <= 1'h0;
      write_done_data_log_force[1758] <= 1'h0;
      write_done_data_log_force[1759] <= 1'h0;
      write_done_data_log_force[1760] <= 1'h0;
      write_done_data_log_force[1761] <= 1'h0;
      write_done_data_log_force[1762] <= 1'h0;
      write_done_data_log_force[1763] <= 1'h0;
      write_done_data_log_force[1764] <= 1'h0;
      write_done_data_log_force[1765] <= 1'h0;
      write_done_data_log_force[1766] <= 1'h0;
      write_done_data_log_force[1767] <= 1'h0;
      write_done_data_log_force[1768] <= 1'h0;
      write_done_data_log_force[1769] <= 1'h0;
      write_done_data_log_force[1770] <= 1'h0;
      write_done_data_log_force[1771] <= 1'h0;
      write_done_data_log_force[1772] <= 1'h0;
      write_done_data_log_force[1773] <= 1'h0;
      write_done_data_log_force[1774] <= 1'h0;
      write_done_data_log_force[1775] <= 1'h0;
      write_done_data_log_force[1776] <= 1'h0;
      write_done_data_log_force[1777] <= 1'h0;
      write_done_data_log_force[1778] <= 1'h0;
      write_done_data_log_force[1779] <= 1'h0;
      write_done_data_log_force[1780] <= 1'h0;
      write_done_data_log_force[1781] <= 1'h0;
      write_done_data_log_force[1782] <= 1'h0;
      write_done_data_log_force[1783] <= 1'h0;
      write_done_data_log_force[1784] <= 1'h0;
      write_done_data_log_force[1785] <= 1'h0;
      write_done_data_log_force[1786] <= 1'h0;
      write_done_data_log_force[1787] <= 1'h0;
      write_done_data_log_force[1788] <= 1'h0;
      write_done_data_log_force[1789] <= 1'h0;
      write_done_data_log_force[1790] <= 1'h0;
      write_done_data_log_force[1791] <= 1'h0;
      write_done_data_log_force[1792] <= 1'h0;
      write_done_data_log_force[1793] <= 1'h0;
      write_done_data_log_force[1794] <= 1'h0;
      write_done_data_log_force[1795] <= 1'h0;
      write_done_data_log_force[1796] <= 1'h0;
      write_done_data_log_force[1797] <= 1'h0;
      write_done_data_log_force[1798] <= 1'h0;
      write_done_data_log_force[1799] <= 1'h0;
      write_done_data_log_force[1800] <= 1'h0;
      write_done_data_log_force[1801] <= 1'h0;
      write_done_data_log_force[1802] <= 1'h0;
      write_done_data_log_force[1803] <= 1'h0;
      write_done_data_log_force[1804] <= 1'h0;
      write_done_data_log_force[1805] <= 1'h0;
      write_done_data_log_force[1806] <= 1'h0;
      write_done_data_log_force[1807] <= 1'h0;
      write_done_data_log_force[1808] <= 1'h0;
      write_done_data_log_force[1809] <= 1'h0;
      write_done_data_log_force[1810] <= 1'h0;
      write_done_data_log_force[1811] <= 1'h0;
      write_done_data_log_force[1812] <= 1'h0;
      write_done_data_log_force[1813] <= 1'h0;
      write_done_data_log_force[1814] <= 1'h0;
      write_done_data_log_force[1815] <= 1'h0;
      write_done_data_log_force[1816] <= 1'h0;
      write_done_data_log_force[1817] <= 1'h0;
      write_done_data_log_force[1818] <= 1'h0;
      write_done_data_log_force[1819] <= 1'h0;
      write_done_data_log_force[1820] <= 1'h0;
      write_done_data_log_force[1821] <= 1'h0;
      write_done_data_log_force[1822] <= 1'h0;
      write_done_data_log_force[1823] <= 1'h0;
      write_done_data_log_force[1824] <= 1'h0;
      write_done_data_log_force[1825] <= 1'h0;
      write_done_data_log_force[1826] <= 1'h0;
      write_done_data_log_force[1827] <= 1'h0;
      write_done_data_log_force[1828] <= 1'h0;
      write_done_data_log_force[1829] <= 1'h0;
      write_done_data_log_force[1830] <= 1'h0;
      write_done_data_log_force[1831] <= 1'h0;
      write_done_data_log_force[1832] <= 1'h0;
      write_done_data_log_force[1833] <= 1'h0;
      write_done_data_log_force[1834] <= 1'h0;
      write_done_data_log_force[1835] <= 1'h0;
      write_done_data_log_force[1836] <= 1'h0;
      write_done_data_log_force[1837] <= 1'h0;
      write_done_data_log_force[1838] <= 1'h0;
      write_done_data_log_force[1839] <= 1'h0;
      write_done_data_log_force[1840] <= 1'h0;
      write_done_data_log_force[1841] <= 1'h0;
      write_done_data_log_force[1842] <= 1'h0;
      write_done_data_log_force[1843] <= 1'h0;
      write_done_data_log_force[1844] <= 1'h0;
      write_done_data_log_force[1845] <= 1'h0;
      write_done_data_log_force[1846] <= 1'h0;
      write_done_data_log_force[1847] <= 1'h0;
      write_done_data_log_force[1848] <= 1'h0;
      write_done_data_log_force[1849] <= 1'h0;
      write_done_data_log_force[1850] <= 1'h0;
      write_done_data_log_force[1851] <= 1'h0;
      write_done_data_log_force[1852] <= 1'h0;
      write_done_data_log_force[1853] <= 1'h0;
      write_done_data_log_force[1854] <= 1'h0;
      write_done_data_log_force[1855] <= 1'h0;
      write_done_data_log_force[1856] <= 1'h0;
      write_done_data_log_force[1857] <= 1'h0;
      write_done_data_log_force[1858] <= 1'h0;
      write_done_data_log_force[1859] <= 1'h0;
      write_done_data_log_force[1860] <= 1'h0;
      write_done_data_log_force[1861] <= 1'h0;
      write_done_data_log_force[1862] <= 1'h0;
      write_done_data_log_force[1863] <= 1'h0;
      write_done_data_log_force[1864] <= 1'h0;
      write_done_data_log_force[1865] <= 1'h0;
      write_done_data_log_force[1866] <= 1'h0;
      write_done_data_log_force[1867] <= 1'h0;
      write_done_data_log_force[1868] <= 1'h0;
      write_done_data_log_force[1869] <= 1'h0;
      write_done_data_log_force[1870] <= 1'h0;
      write_done_data_log_force[1871] <= 1'h0;
      write_done_data_log_force[1872] <= 1'h0;
      write_done_data_log_force[1873] <= 1'h0;
      write_done_data_log_force[1874] <= 1'h0;
      write_done_data_log_force[1875] <= 1'h0;
      write_done_data_log_force[1876] <= 1'h0;
      write_done_data_log_force[1877] <= 1'h0;
      write_done_data_log_force[1878] <= 1'h0;
      write_done_data_log_force[1879] <= 1'h0;
      write_done_data_log_force[1880] <= 1'h0;
      write_done_data_log_force[1881] <= 1'h0;
      write_done_data_log_force[1882] <= 1'h0;
      write_done_data_log_force[1883] <= 1'h0;
      write_done_data_log_force[1884] <= 1'h0;
      write_done_data_log_force[1885] <= 1'h0;
      write_done_data_log_force[1886] <= 1'h0;
      write_done_data_log_force[1887] <= 1'h0;
      write_done_data_log_force[1888] <= 1'h0;
      write_done_data_log_force[1889] <= 1'h0;
      write_done_data_log_force[1890] <= 1'h0;
      write_done_data_log_force[1891] <= 1'h0;
      write_done_data_log_force[1892] <= 1'h0;
      write_done_data_log_force[1893] <= 1'h0;
      write_done_data_log_force[1894] <= 1'h0;
      write_done_data_log_force[1895] <= 1'h0;
      write_done_data_log_force[1896] <= 1'h0;
      write_done_data_log_force[1897] <= 1'h0;
      write_done_data_log_force[1898] <= 1'h0;
      write_done_data_log_force[1899] <= 1'h0;
      write_done_data_log_force[1900] <= 1'h0;
      write_done_data_log_force[1901] <= 1'h0;
      write_done_data_log_force[1902] <= 1'h0;
      write_done_data_log_force[1903] <= 1'h0;
      write_done_data_log_force[1904] <= 1'h0;
      write_done_data_log_force[1905] <= 1'h0;
      write_done_data_log_force[1906] <= 1'h0;
      write_done_data_log_force[1907] <= 1'h0;
      write_done_data_log_force[1908] <= 1'h0;
      write_done_data_log_force[1909] <= 1'h0;
      write_done_data_log_force[1910] <= 1'h0;
      write_done_data_log_force[1911] <= 1'h0;
      write_done_data_log_force[1912] <= 1'h0;
      write_done_data_log_force[1913] <= 1'h0;
      write_done_data_log_force[1914] <= 1'h0;
      write_done_data_log_force[1915] <= 1'h0;
      write_done_data_log_force[1916] <= 1'h0;
      write_done_data_log_force[1917] <= 1'h0;
      write_done_data_log_force[1918] <= 1'h0;
      write_done_data_log_force[1919] <= 1'h0;
      write_done_data_log_force[1920] <= 1'h0;
      write_done_data_log_force[1921] <= 1'h0;
      write_done_data_log_force[1922] <= 1'h0;
      write_done_data_log_force[1923] <= 1'h0;
      write_done_data_log_force[1924] <= 1'h0;
      write_done_data_log_force[1925] <= 1'h0;
      write_done_data_log_force[1926] <= 1'h0;
      write_done_data_log_force[1927] <= 1'h0;
      write_done_data_log_force[1928] <= 1'h0;
      write_done_data_log_force[1929] <= 1'h0;
      write_done_data_log_force[1930] <= 1'h0;
      write_done_data_log_force[1931] <= 1'h0;
      write_done_data_log_force[1932] <= 1'h0;
      write_done_data_log_force[1933] <= 1'h0;
      write_done_data_log_force[1934] <= 1'h0;
      write_done_data_log_force[1935] <= 1'h0;
      write_done_data_log_force[1936] <= 1'h0;
      write_done_data_log_force[1937] <= 1'h0;
      write_done_data_log_force[1938] <= 1'h0;
      write_done_data_log_force[1939] <= 1'h0;
      write_done_data_log_force[1940] <= 1'h0;
      write_done_data_log_force[1941] <= 1'h0;
      write_done_data_log_force[1942] <= 1'h0;
      write_done_data_log_force[1943] <= 1'h0;
      write_done_data_log_force[1944] <= 1'h0;
      write_done_data_log_force[1945] <= 1'h0;
      write_done_data_log_force[1946] <= 1'h0;
      write_done_data_log_force[1947] <= 1'h0;
      write_done_data_log_force[1948] <= 1'h0;
      write_done_data_log_force[1949] <= 1'h0;
      write_done_data_log_force[1950] <= 1'h0;
      write_done_data_log_force[1951] <= 1'h0;
      write_done_data_log_force[1952] <= 1'h0;
      write_done_data_log_force[1953] <= 1'h0;
      write_done_data_log_force[1954] <= 1'h0;
      write_done_data_log_force[1955] <= 1'h0;
      write_done_data_log_force[1956] <= 1'h0;
      write_done_data_log_force[1957] <= 1'h0;
      write_done_data_log_force[1958] <= 1'h0;
      write_done_data_log_force[1959] <= 1'h0;
      write_done_data_log_force[1960] <= 1'h0;
      write_done_data_log_force[1961] <= 1'h0;
      write_done_data_log_force[1962] <= 1'h0;
      write_done_data_log_force[1963] <= 1'h0;
      write_done_data_log_force[1964] <= 1'h0;
      write_done_data_log_force[1965] <= 1'h0;
      write_done_data_log_force[1966] <= 1'h0;
      write_done_data_log_force[1967] <= 1'h0;
      write_done_data_log_force[1968] <= 1'h0;
      write_done_data_log_force[1969] <= 1'h0;
      write_done_data_log_force[1970] <= 1'h0;
      write_done_data_log_force[1971] <= 1'h0;
      write_done_data_log_force[1972] <= 1'h0;
      write_done_data_log_force[1973] <= 1'h0;
      write_done_data_log_force[1974] <= 1'h0;
      write_done_data_log_force[1975] <= 1'h0;
      write_done_data_log_force[1976] <= 1'h0;
      write_done_data_log_force[1977] <= 1'h0;
      write_done_data_log_force[1978] <= 1'h0;
      write_done_data_log_force[1979] <= 1'h0;
      write_done_data_log_force[1980] <= 1'h0;
      write_done_data_log_force[1981] <= 1'h0;
      write_done_data_log_force[1982] <= 1'h0;
      write_done_data_log_force[1983] <= 1'h0;
      write_done_data_log_force[1984] <= 1'h0;
      write_done_data_log_force[1985] <= 1'h0;
      write_done_data_log_force[1986] <= 1'h0;
      write_done_data_log_force[1987] <= 1'h0;
      write_done_data_log_force[1988] <= 1'h0;
      write_done_data_log_force[1989] <= 1'h0;
      write_done_data_log_force[1990] <= 1'h0;
      write_done_data_log_force[1991] <= 1'h0;
      write_done_data_log_force[1992] <= 1'h0;
      write_done_data_log_force[1993] <= 1'h0;
      write_done_data_log_force[1994] <= 1'h0;
      write_done_data_log_force[1995] <= 1'h0;
      write_done_data_log_force[1996] <= 1'h0;
      write_done_data_log_force[1997] <= 1'h0;
      write_done_data_log_force[1998] <= 1'h0;
      write_done_data_log_force[1999] <= 1'h0;
      write_done_data_log_force[2000] <= 1'h0;
      write_done_data_log_force[2001] <= 1'h0;
      write_done_data_log_force[2002] <= 1'h0;
      write_done_data_log_force[2003] <= 1'h0;
      write_done_data_log_force[2004] <= 1'h0;
      write_done_data_log_force[2005] <= 1'h0;
      write_done_data_log_force[2006] <= 1'h0;
      write_done_data_log_force[2007] <= 1'h0;
      write_done_data_log_force[2008] <= 1'h0;
      write_done_data_log_force[2009] <= 1'h0;
      write_done_data_log_force[2010] <= 1'h0;
      write_done_data_log_force[2011] <= 1'h0;
      write_done_data_log_force[2012] <= 1'h0;
      write_done_data_log_force[2013] <= 1'h0;
      write_done_data_log_force[2014] <= 1'h0;
      write_done_data_log_force[2015] <= 1'h0;
      write_done_data_log_force[2016] <= 1'h0;
      write_done_data_log_force[2017] <= 1'h0;
      write_done_data_log_force[2018] <= 1'h0;
      write_done_data_log_force[2019] <= 1'h0;
      write_done_data_log_force[2020] <= 1'h0;
      write_done_data_log_force[2021] <= 1'h0;
      write_done_data_log_force[2022] <= 1'h0;
      write_done_data_log_force[2023] <= 1'h0;
      write_done_data_log_force[2024] <= 1'h0;
      write_done_data_log_force[2025] <= 1'h0;
      write_done_data_log_force[2026] <= 1'h0;
      write_done_data_log_force[2027] <= 1'h0;
      write_done_data_log_force[2028] <= 1'h0;
      write_done_data_log_force[2029] <= 1'h0;
      write_done_data_log_force[2030] <= 1'h0;
      write_done_data_log_force[2031] <= 1'h0;
      write_done_data_log_force[2032] <= 1'h0;
      write_done_data_log_force[2033] <= 1'h0;
      write_done_data_log_force[2034] <= 1'h0;
      write_done_data_log_force[2035] <= 1'h0;
      write_done_data_log_force[2036] <= 1'h0;
      write_done_data_log_force[2037] <= 1'h0;
      write_done_data_log_force[2038] <= 1'h0;
      write_done_data_log_force[2039] <= 1'h0;
      write_done_data_log_force[2040] <= 1'h0;
      write_done_data_log_force[2041] <= 1'h0;
      write_done_data_log_force[2042] <= 1'h0;
      write_done_data_log_force[2043] <= 1'h0;
      write_done_data_log_force[2044] <= 1'h0;
      write_done_data_log_force[2045] <= 1'h0;
      write_done_data_log_force[2046] <= 1'h0;
      write_done_data_log_force[2047] <= 1'h0;
      write_done_data_log_force[2048] <= 1'h0;
      write_done_data_log_force[2049] <= 1'h0;
      write_done_data_log_force[2050] <= 1'h0;
      write_done_data_log_force[2051] <= 1'h0;
      write_done_data_log_force[2052] <= 1'h0;
      write_done_data_log_force[2053] <= 1'h0;
      write_done_data_log_force[2054] <= 1'h0;
      write_done_data_log_force[2055] <= 1'h0;
      write_done_data_log_force[2056] <= 1'h0;
      write_done_data_log_force[2057] <= 1'h0;
      write_done_data_log_force[2058] <= 1'h0;
      write_done_data_log_force[2059] <= 1'h0;
      write_done_data_log_force[2060] <= 1'h0;
      write_done_data_log_force[2061] <= 1'h0;
      write_done_data_log_force[2062] <= 1'h0;
      write_done_data_log_force[2063] <= 1'h0;
      write_done_data_log_force[2064] <= 1'h0;
      write_done_data_log_force[2065] <= 1'h0;
      write_done_data_log_force[2066] <= 1'h0;
      write_done_data_log_force[2067] <= 1'h0;
      write_done_data_log_force[2068] <= 1'h0;
      write_done_data_log_force[2069] <= 1'h0;
      write_done_data_log_force[2070] <= 1'h0;
      write_done_data_log_force[2071] <= 1'h0;
      write_done_data_log_force[2072] <= 1'h0;
      write_done_data_log_force[2073] <= 1'h0;
      write_done_data_log_force[2074] <= 1'h0;
      write_done_data_log_force[2075] <= 1'h0;
      write_done_data_log_force[2076] <= 1'h0;
      write_done_data_log_force[2077] <= 1'h0;
      write_done_data_log_force[2078] <= 1'h0;
      write_done_data_log_force[2079] <= 1'h0;
      write_done_data_log_force[2080] <= 1'h0;
      write_done_data_log_force[2081] <= 1'h0;
      write_done_data_log_force[2082] <= 1'h0;
      write_done_data_log_force[2083] <= 1'h0;
      write_done_data_log_force[2084] <= 1'h0;
      write_done_data_log_force[2085] <= 1'h0;
      write_done_data_log_force[2086] <= 1'h0;
      write_done_data_log_force[2087] <= 1'h0;
      write_done_data_log_force[2088] <= 1'h0;
      write_done_data_log_force[2089] <= 1'h0;
      write_done_data_log_force[2090] <= 1'h0;
      write_done_data_log_force[2091] <= 1'h0;
      write_done_data_log_force[2092] <= 1'h0;
      write_done_data_log_force[2093] <= 1'h0;
      write_done_data_log_force[2094] <= 1'h0;
      write_done_data_log_force[2095] <= 1'h0;
      write_done_data_log_force[2096] <= 1'h0;
      write_done_data_log_force[2097] <= 1'h0;
      write_done_data_log_force[2098] <= 1'h0;
      write_done_data_log_force[2099] <= 1'h0;
      write_done_data_log_force[2100] <= 1'h0;
      write_done_data_log_force[2101] <= 1'h0;
      write_done_data_log_force[2102] <= 1'h0;
      write_done_data_log_force[2103] <= 1'h0;
      write_done_data_log_force[2104] <= 1'h0;
      write_done_data_log_force[2105] <= 1'h0;
      write_done_data_log_force[2106] <= 1'h0;
      write_done_data_log_force[2107] <= 1'h0;
      write_done_data_log_force[2108] <= 1'h0;
      write_done_data_log_force[2109] <= 1'h0;
      write_done_data_log_force[2110] <= 1'h0;
      write_done_data_log_force[2111] <= 1'h0;
      write_done_data_log_force[2112] <= 1'h0;
      write_done_data_log_force[2113] <= 1'h0;
      write_done_data_log_force[2114] <= 1'h0;
      write_done_data_log_force[2115] <= 1'h0;
      write_done_data_log_force[2116] <= 1'h0;
      write_done_data_log_force[2117] <= 1'h0;
      write_done_data_log_force[2118] <= 1'h0;
      write_done_data_log_force[2119] <= 1'h0;
      write_done_data_log_force[2120] <= 1'h0;
      write_done_data_log_force[2121] <= 1'h0;
      write_done_data_log_force[2122] <= 1'h0;
      write_done_data_log_force[2123] <= 1'h0;
      write_done_data_log_force[2124] <= 1'h0;
      write_done_data_log_force[2125] <= 1'h0;
      write_done_data_log_force[2126] <= 1'h0;
      write_done_data_log_force[2127] <= 1'h0;
      write_done_data_log_force[2128] <= 1'h0;
      write_done_data_log_force[2129] <= 1'h0;
      write_done_data_log_force[2130] <= 1'h0;
      write_done_data_log_force[2131] <= 1'h0;
      write_done_data_log_force[2132] <= 1'h0;
      write_done_data_log_force[2133] <= 1'h0;
      write_done_data_log_force[2134] <= 1'h0;
      write_done_data_log_force[2135] <= 1'h0;
      write_done_data_log_force[2136] <= 1'h0;
      write_done_data_log_force[2137] <= 1'h0;
      write_done_data_log_force[2138] <= 1'h0;
      write_done_data_log_force[2139] <= 1'h0;
      write_done_data_log_force[2140] <= 1'h0;
      write_done_data_log_force[2141] <= 1'h0;
      write_done_data_log_force[2142] <= 1'h0;
      write_done_data_log_force[2143] <= 1'h0;
      write_done_data_log_force[2144] <= 1'h0;
      write_done_data_log_force[2145] <= 1'h0;
      write_done_data_log_force[2146] <= 1'h0;
      write_done_data_log_force[2147] <= 1'h0;
      write_done_data_log_force[2148] <= 1'h0;
      write_done_data_log_force[2149] <= 1'h0;
      write_done_data_log_force[2150] <= 1'h0;
      write_done_data_log_force[2151] <= 1'h0;
      write_done_data_log_force[2152] <= 1'h0;
      write_done_data_log_force[2153] <= 1'h0;
      write_done_data_log_force[2154] <= 1'h0;
      write_done_data_log_force[2155] <= 1'h0;
      write_done_data_log_force[2156] <= 1'h0;
      write_done_data_log_force[2157] <= 1'h0;
      write_done_data_log_force[2158] <= 1'h0;
      write_done_data_log_force[2159] <= 1'h0;
      write_done_data_log_force[2160] <= 1'h0;
      write_done_data_log_force[2161] <= 1'h0;
      write_done_data_log_force[2162] <= 1'h0;
      write_done_data_log_force[2163] <= 1'h0;
      write_done_data_log_force[2164] <= 1'h0;
      write_done_data_log_force[2165] <= 1'h0;
      write_done_data_log_force[2166] <= 1'h0;
      write_done_data_log_force[2167] <= 1'h0;
      write_done_data_log_force[2168] <= 1'h0;
      write_done_data_log_force[2169] <= 1'h0;
      write_done_data_log_force[2170] <= 1'h0;
      write_done_data_log_force[2171] <= 1'h0;
      write_done_data_log_force[2172] <= 1'h0;
      write_done_data_log_force[2173] <= 1'h0;
      write_done_data_log_force[2174] <= 1'h0;
      write_done_data_log_force[2175] <= 1'h0;
      write_done_data_log_force[2176] <= 1'h0;
      write_done_data_log_force[2177] <= 1'h0;
      write_done_data_log_force[2178] <= 1'h0;
      write_done_data_log_force[2179] <= 1'h0;
      write_done_data_log_force[2180] <= 1'h0;
      write_done_data_log_force[2181] <= 1'h0;
      write_done_data_log_force[2182] <= 1'h0;
      write_done_data_log_force[2183] <= 1'h0;
      write_done_data_log_force[2184] <= 1'h0;
      write_done_data_log_force[2185] <= 1'h0;
      write_done_data_log_force[2186] <= 1'h0;
      write_done_data_log_force[2187] <= 1'h0;
      write_done_data_log_force[2188] <= 1'h0;
      write_done_data_log_force[2189] <= 1'h0;
      write_done_data_log_force[2190] <= 1'h0;
      write_done_data_log_force[2191] <= 1'h0;
      write_done_data_log_force[2192] <= 1'h0;
      write_done_data_log_force[2193] <= 1'h0;
      write_done_data_log_force[2194] <= 1'h0;
      write_done_data_log_force[2195] <= 1'h0;
      write_done_data_log_force[2196] <= 1'h0;
      write_done_data_log_force[2197] <= 1'h0;
      write_done_data_log_force[2198] <= 1'h0;
      write_done_data_log_force[2199] <= 1'h0;
      write_done_data_log_force[2200] <= 1'h0;
      write_done_data_log_force[2201] <= 1'h0;
      write_done_data_log_force[2202] <= 1'h0;
      write_done_data_log_force[2203] <= 1'h0;
      write_done_data_log_force[2204] <= 1'h0;
      write_done_data_log_force[2205] <= 1'h0;
      write_done_data_log_force[2206] <= 1'h0;
      write_done_data_log_force[2207] <= 1'h0;
      write_done_data_log_force[2208] <= 1'h0;
      write_done_data_log_force[2209] <= 1'h0;
      write_done_data_log_force[2210] <= 1'h0;
      write_done_data_log_force[2211] <= 1'h0;
      write_done_data_log_force[2212] <= 1'h0;
      write_done_data_log_force[2213] <= 1'h0;
      write_done_data_log_force[2214] <= 1'h0;
      write_done_data_log_force[2215] <= 1'h0;
      write_done_data_log_force[2216] <= 1'h0;
      write_done_data_log_force[2217] <= 1'h0;
      write_done_data_log_force[2218] <= 1'h0;
      write_done_data_log_force[2219] <= 1'h0;
      write_done_data_log_force[2220] <= 1'h0;
      write_done_data_log_force[2221] <= 1'h0;
      write_done_data_log_force[2222] <= 1'h0;
      write_done_data_log_force[2223] <= 1'h0;
      write_done_data_log_force[2224] <= 1'h0;
      write_done_data_log_force[2225] <= 1'h0;
      write_done_data_log_force[2226] <= 1'h0;
      write_done_data_log_force[2227] <= 1'h0;
      write_done_data_log_force[2228] <= 1'h0;
      write_done_data_log_force[2229] <= 1'h0;
      write_done_data_log_force[2230] <= 1'h0;
      write_done_data_log_force[2231] <= 1'h0;
      write_done_data_log_force[2232] <= 1'h0;
      write_done_data_log_force[2233] <= 1'h0;
      write_done_data_log_force[2234] <= 1'h0;
      write_done_data_log_force[2235] <= 1'h0;
      write_done_data_log_force[2236] <= 1'h0;
      write_done_data_log_force[2237] <= 1'h0;
      write_done_data_log_force[2238] <= 1'h0;
      write_done_data_log_force[2239] <= 1'h0;
      write_done_data_log_force[2240] <= 1'h0;
      write_done_data_log_force[2241] <= 1'h0;
      write_done_data_log_force[2242] <= 1'h0;
      write_done_data_log_force[2243] <= 1'h0;
      write_done_data_log_force[2244] <= 1'h0;
      write_done_data_log_force[2245] <= 1'h0;
      write_done_data_log_force[2246] <= 1'h0;
      write_done_data_log_force[2247] <= 1'h0;
      write_done_data_log_force[2248] <= 1'h0;
      write_done_data_log_force[2249] <= 1'h0;
      write_done_data_log_force[2250] <= 1'h0;
      write_done_data_log_force[2251] <= 1'h0;
      write_done_data_log_force[2252] <= 1'h0;
      write_done_data_log_force[2253] <= 1'h0;
      write_done_data_log_force[2254] <= 1'h0;
      write_done_data_log_force[2255] <= 1'h0;
      write_done_data_log_force[2256] <= 1'h0;
      write_done_data_log_force[2257] <= 1'h0;
      write_done_data_log_force[2258] <= 1'h0;
      write_done_data_log_force[2259] <= 1'h0;
      write_done_data_log_force[2260] <= 1'h0;
      write_done_data_log_force[2261] <= 1'h0;
      write_done_data_log_force[2262] <= 1'h0;
      write_done_data_log_force[2263] <= 1'h0;
      write_done_data_log_force[2264] <= 1'h0;
      write_done_data_log_force[2265] <= 1'h0;
      write_done_data_log_force[2266] <= 1'h0;
      write_done_data_log_force[2267] <= 1'h0;
      write_done_data_log_force[2268] <= 1'h0;
      write_done_data_log_force[2269] <= 1'h0;
      write_done_data_log_force[2270] <= 1'h0;
      write_done_data_log_force[2271] <= 1'h0;
      write_done_data_log_force[2272] <= 1'h0;
      write_done_data_log_force[2273] <= 1'h0;
      write_done_data_log_force[2274] <= 1'h0;
      write_done_data_log_force[2275] <= 1'h0;
      write_done_data_log_force[2276] <= 1'h0;
      write_done_data_log_force[2277] <= 1'h0;
      write_done_data_log_force[2278] <= 1'h0;
      write_done_data_log_force[2279] <= 1'h0;
      write_done_data_log_force[2280] <= 1'h0;
      write_done_data_log_force[2281] <= 1'h0;
      write_done_data_log_force[2282] <= 1'h0;
      write_done_data_log_force[2283] <= 1'h0;
      write_done_data_log_force[2284] <= 1'h0;
      write_done_data_log_force[2285] <= 1'h0;
      write_done_data_log_force[2286] <= 1'h0;
      write_done_data_log_force[2287] <= 1'h0;
      write_done_data_log_force[2288] <= 1'h0;
      write_done_data_log_force[2289] <= 1'h0;
      write_done_data_log_force[2290] <= 1'h0;
      write_done_data_log_force[2291] <= 1'h0;
      write_done_data_log_force[2292] <= 1'h0;
      write_done_data_log_force[2293] <= 1'h0;
      write_done_data_log_force[2294] <= 1'h0;
      write_done_data_log_force[2295] <= 1'h0;
      write_done_data_log_force[2296] <= 1'h0;
      write_done_data_log_force[2297] <= 1'h0;
      write_done_data_log_force[2298] <= 1'h0;
      write_done_data_log_force[2299] <= 1'h0;
      write_done_data_log_force[2300] <= 1'h0;
      write_done_data_log_force[2301] <= 1'h0;
      write_done_data_log_force[2302] <= 1'h0;
      write_done_data_log_force[2303] <= 1'h0;
      write_done_data_log_force[2304] <= 1'h0;
      write_done_data_log_force[2305] <= 1'h0;
      write_done_data_log_force[2306] <= 1'h0;
      write_done_data_log_force[2307] <= 1'h0;
      write_done_data_log_force[2308] <= 1'h0;
      write_done_data_log_force[2309] <= 1'h0;
      write_done_data_log_force[2310] <= 1'h0;
      write_done_data_log_force[2311] <= 1'h0;
      write_done_data_log_force[2312] <= 1'h0;
      write_done_data_log_force[2313] <= 1'h0;
      write_done_data_log_force[2314] <= 1'h0;
      write_done_data_log_force[2315] <= 1'h0;
      write_done_data_log_force[2316] <= 1'h0;
      write_done_data_log_force[2317] <= 1'h0;
      write_done_data_log_force[2318] <= 1'h0;
      write_done_data_log_force[2319] <= 1'h0;
      write_done_data_log_force[2320] <= 1'h0;
      write_done_data_log_force[2321] <= 1'h0;
      write_done_data_log_force[2322] <= 1'h0;
      write_done_data_log_force[2323] <= 1'h0;
      write_done_data_log_force[2324] <= 1'h0;
      write_done_data_log_force[2325] <= 1'h0;
      write_done_data_log_force[2326] <= 1'h0;
      write_done_data_log_force[2327] <= 1'h0;
      write_done_data_log_force[2328] <= 1'h0;
      write_done_data_log_force[2329] <= 1'h0;
      write_done_data_log_force[2330] <= 1'h0;
      write_done_data_log_force[2331] <= 1'h0;
      write_done_data_log_force[2332] <= 1'h0;
      write_done_data_log_force[2333] <= 1'h0;
      write_done_data_log_force[2334] <= 1'h0;
      write_done_data_log_force[2335] <= 1'h0;
      write_done_data_log_force[2336] <= 1'h0;
      write_done_data_log_force[2337] <= 1'h0;
      write_done_data_log_force[2338] <= 1'h0;
      write_done_data_log_force[2339] <= 1'h0;
      write_done_data_log_force[2340] <= 1'h0;
      write_done_data_log_force[2341] <= 1'h0;
      write_done_data_log_force[2342] <= 1'h0;
      write_done_data_log_force[2343] <= 1'h0;
      write_done_data_log_force[2344] <= 1'h0;
      write_done_data_log_force[2345] <= 1'h0;
      write_done_data_log_force[2346] <= 1'h0;
      write_done_data_log_force[2347] <= 1'h0;
      write_done_data_log_force[2348] <= 1'h0;
      write_done_data_log_force[2349] <= 1'h0;
      write_done_data_log_force[2350] <= 1'h0;
      write_done_data_log_force[2351] <= 1'h0;
      write_done_data_log_force[2352] <= 1'h0;
      write_done_data_log_force[2353] <= 1'h0;
      write_done_data_log_force[2354] <= 1'h0;
      write_done_data_log_force[2355] <= 1'h0;
      write_done_data_log_force[2356] <= 1'h0;
      write_done_data_log_force[2357] <= 1'h0;
      write_done_data_log_force[2358] <= 1'h0;
      write_done_data_log_force[2359] <= 1'h0;
      write_done_data_log_force[2360] <= 1'h0;
      write_done_data_log_force[2361] <= 1'h0;
      write_done_data_log_force[2362] <= 1'h0;
      write_done_data_log_force[2363] <= 1'h0;
      write_done_data_log_force[2364] <= 1'h0;
      write_done_data_log_force[2365] <= 1'h0;
      write_done_data_log_force[2366] <= 1'h0;
      write_done_data_log_force[2367] <= 1'h0;
      write_done_data_log_force[2368] <= 1'h0;
      write_done_data_log_force[2369] <= 1'h0;
      write_done_data_log_force[2370] <= 1'h0;
      write_done_data_log_force[2371] <= 1'h0;
      write_done_data_log_force[2372] <= 1'h0;
      write_done_data_log_force[2373] <= 1'h0;
      write_done_data_log_force[2374] <= 1'h0;
      write_done_data_log_force[2375] <= 1'h0;
      write_done_data_log_force[2376] <= 1'h0;
      write_done_data_log_force[2377] <= 1'h0;
      write_done_data_log_force[2378] <= 1'h0;
      write_done_data_log_force[2379] <= 1'h0;
      write_done_data_log_force[2380] <= 1'h0;
      write_done_data_log_force[2381] <= 1'h0;
      write_done_data_log_force[2382] <= 1'h0;
      write_done_data_log_force[2383] <= 1'h0;
      write_done_data_log_force[2384] <= 1'h0;
      write_done_data_log_force[2385] <= 1'h0;
      write_done_data_log_force[2386] <= 1'h0;
      write_done_data_log_force[2387] <= 1'h0;
      write_done_data_log_force[2388] <= 1'h0;
      write_done_data_log_force[2389] <= 1'h0;
      write_done_data_log_force[2390] <= 1'h0;
      write_done_data_log_force[2391] <= 1'h0;
      write_done_data_log_force[2392] <= 1'h0;
      write_done_data_log_force[2393] <= 1'h0;
      write_done_data_log_force[2394] <= 1'h0;
      write_done_data_log_force[2395] <= 1'h0;
      write_done_data_log_force[2396] <= 1'h0;
      write_done_data_log_force[2397] <= 1'h0;
      write_done_data_log_force[2398] <= 1'h0;
      write_done_data_log_force[2399] <= 1'h0;
      write_done_data_log_force[2400] <= 1'h0;
      write_done_data_log_force[2401] <= 1'h0;
      write_done_data_log_force[2402] <= 1'h0;
      write_done_data_log_force[2403] <= 1'h0;
      write_done_data_log_force[2404] <= 1'h0;
      write_done_data_log_force[2405] <= 1'h0;
      write_done_data_log_force[2406] <= 1'h0;
      write_done_data_log_force[2407] <= 1'h0;
      write_done_data_log_force[2408] <= 1'h0;
      write_done_data_log_force[2409] <= 1'h0;
      write_done_data_log_force[2410] <= 1'h0;
      write_done_data_log_force[2411] <= 1'h0;
      write_done_data_log_force[2412] <= 1'h0;
      write_done_data_log_force[2413] <= 1'h0;
      write_done_data_log_force[2414] <= 1'h0;
      write_done_data_log_force[2415] <= 1'h0;
      write_done_data_log_force[2416] <= 1'h0;
      write_done_data_log_force[2417] <= 1'h0;
      write_done_data_log_force[2418] <= 1'h0;
      write_done_data_log_force[2419] <= 1'h0;
      write_done_data_log_force[2420] <= 1'h0;
      write_done_data_log_force[2421] <= 1'h0;
      write_done_data_log_force[2422] <= 1'h0;
      write_done_data_log_force[2423] <= 1'h0;
      write_done_data_log_force[2424] <= 1'h0;
      write_done_data_log_force[2425] <= 1'h0;
      write_done_data_log_force[2426] <= 1'h0;
      write_done_data_log_force[2427] <= 1'h0;
      write_done_data_log_force[2428] <= 1'h0;
      write_done_data_log_force[2429] <= 1'h0;
      write_done_data_log_force[2430] <= 1'h0;
      write_done_data_log_force[2431] <= 1'h0;
      write_done_data_log_force[2432] <= 1'h0;
      write_done_data_log_force[2433] <= 1'h0;
      write_done_data_log_force[2434] <= 1'h0;
      write_done_data_log_force[2435] <= 1'h0;
      write_done_data_log_force[2436] <= 1'h0;
      write_done_data_log_force[2437] <= 1'h0;
      write_done_data_log_force[2438] <= 1'h0;
      write_done_data_log_force[2439] <= 1'h0;
      write_done_data_log_force[2440] <= 1'h0;
      write_done_data_log_force[2441] <= 1'h0;
      write_done_data_log_force[2442] <= 1'h0;
      write_done_data_log_force[2443] <= 1'h0;
      write_done_data_log_force[2444] <= 1'h0;
      write_done_data_log_force[2445] <= 1'h0;
      write_done_data_log_force[2446] <= 1'h0;
      write_done_data_log_force[2447] <= 1'h0;
      write_done_data_log_force[2448] <= 1'h0;
      write_done_data_log_force[2449] <= 1'h0;
      write_done_data_log_force[2450] <= 1'h0;
      write_done_data_log_force[2451] <= 1'h0;
      write_done_data_log_force[2452] <= 1'h0;
      write_done_data_log_force[2453] <= 1'h0;
      write_done_data_log_force[2454] <= 1'h0;
      write_done_data_log_force[2455] <= 1'h0;
      write_done_data_log_force[2456] <= 1'h0;
      write_done_data_log_force[2457] <= 1'h0;
      write_done_data_log_force[2458] <= 1'h0;
      write_done_data_log_force[2459] <= 1'h0;
      write_done_data_log_force[2460] <= 1'h0;
      write_done_data_log_force[2461] <= 1'h0;
      write_done_data_log_force[2462] <= 1'h0;
      write_done_data_log_force[2463] <= 1'h0;
      write_done_data_log_force[2464] <= 1'h0;
      write_done_data_log_force[2465] <= 1'h0;
      write_done_data_log_force[2466] <= 1'h0;
      write_done_data_log_force[2467] <= 1'h0;
      write_done_data_log_force[2468] <= 1'h0;
      write_done_data_log_force[2469] <= 1'h0;
      write_done_data_log_force[2470] <= 1'h0;
      write_done_data_log_force[2471] <= 1'h0;
      write_done_data_log_force[2472] <= 1'h0;
      write_done_data_log_force[2473] <= 1'h0;
      write_done_data_log_force[2474] <= 1'h0;
      write_done_data_log_force[2475] <= 1'h0;
      write_done_data_log_force[2476] <= 1'h0;
      write_done_data_log_force[2477] <= 1'h0;
      write_done_data_log_force[2478] <= 1'h0;
      write_done_data_log_force[2479] <= 1'h0;
      write_done_data_log_force[2480] <= 1'h0;
      write_done_data_log_force[2481] <= 1'h0;
      write_done_data_log_force[2482] <= 1'h0;
      write_done_data_log_force[2483] <= 1'h0;
      write_done_data_log_force[2484] <= 1'h0;
      write_done_data_log_force[2485] <= 1'h0;
      write_done_data_log_force[2486] <= 1'h0;
      write_done_data_log_force[2487] <= 1'h0;
      write_done_data_log_force[2488] <= 1'h0;
      write_done_data_log_force[2489] <= 1'h0;
      write_done_data_log_force[2490] <= 1'h0;
      write_done_data_log_force[2491] <= 1'h0;
      write_done_data_log_force[2492] <= 1'h0;
      write_done_data_log_force[2493] <= 1'h0;
      write_done_data_log_force[2494] <= 1'h0;
      write_done_data_log_force[2495] <= 1'h0;
      write_done_data_log_force[2496] <= 1'h0;
      write_done_data_log_force[2497] <= 1'h0;
      write_done_data_log_force[2498] <= 1'h0;
      write_done_data_log_force[2499] <= 1'h0;
      write_done_data_log_force[2500] <= 1'h0;
      write_done_data_log_force[2501] <= 1'h0;
      write_done_data_log_force[2502] <= 1'h0;
      write_done_data_log_force[2503] <= 1'h0;
      write_done_data_log_force[2504] <= 1'h0;
      write_done_data_log_force[2505] <= 1'h0;
      write_done_data_log_force[2506] <= 1'h0;
      write_done_data_log_force[2507] <= 1'h0;
      write_done_data_log_force[2508] <= 1'h0;
      write_done_data_log_force[2509] <= 1'h0;
      write_done_data_log_force[2510] <= 1'h0;
      write_done_data_log_force[2511] <= 1'h0;
      write_done_data_log_force[2512] <= 1'h0;
      write_done_data_log_force[2513] <= 1'h0;
      write_done_data_log_force[2514] <= 1'h0;
      write_done_data_log_force[2515] <= 1'h0;
      write_done_data_log_force[2516] <= 1'h0;
      write_done_data_log_force[2517] <= 1'h0;
      write_done_data_log_force[2518] <= 1'h0;
      write_done_data_log_force[2519] <= 1'h0;
      write_done_data_log_force[2520] <= 1'h0;
      write_done_data_log_force[2521] <= 1'h0;
      write_done_data_log_force[2522] <= 1'h0;
      write_done_data_log_force[2523] <= 1'h0;
      write_done_data_log_force[2524] <= 1'h0;
      write_done_data_log_force[2525] <= 1'h0;
      write_done_data_log_force[2526] <= 1'h0;
      write_done_data_log_force[2527] <= 1'h0;
      write_done_data_log_force[2528] <= 1'h0;
      write_done_data_log_force[2529] <= 1'h0;
      write_done_data_log_force[2530] <= 1'h0;
      write_done_data_log_force[2531] <= 1'h0;
      write_done_data_log_force[2532] <= 1'h0;
      write_done_data_log_force[2533] <= 1'h0;
      write_done_data_log_force[2534] <= 1'h0;
      write_done_data_log_force[2535] <= 1'h0;
      write_done_data_log_force[2536] <= 1'h0;
      write_done_data_log_force[2537] <= 1'h0;
      write_done_data_log_force[2538] <= 1'h0;
      write_done_data_log_force[2539] <= 1'h0;
      write_done_data_log_force[2540] <= 1'h0;
      write_done_data_log_force[2541] <= 1'h0;
      write_done_data_log_force[2542] <= 1'h0;
      write_done_data_log_force[2543] <= 1'h0;
      write_done_data_log_force[2544] <= 1'h0;
      write_done_data_log_force[2545] <= 1'h0;
      write_done_data_log_force[2546] <= 1'h0;
      write_done_data_log_force[2547] <= 1'h0;
      write_done_data_log_force[2548] <= 1'h0;
      write_done_data_log_force[2549] <= 1'h0;
      write_done_data_log_force[2550] <= 1'h0;
      write_done_data_log_force[2551] <= 1'h0;
      write_done_data_log_force[2552] <= 1'h0;
      write_done_data_log_force[2553] <= 1'h0;
      write_done_data_log_force[2554] <= 1'h0;
      write_done_data_log_force[2555] <= 1'h0;
      write_done_data_log_force[2556] <= 1'h0;
      write_done_data_log_force[2557] <= 1'h0;
      write_done_data_log_force[2558] <= 1'h0;
      write_done_data_log_force[2559] <= 1'h0;
      write_done_data_log_force[2560] <= 1'h0;
      write_done_data_log_force[2561] <= 1'h0;
      write_done_data_log_force[2562] <= 1'h0;
      write_done_data_log_force[2563] <= 1'h0;
      write_done_data_log_force[2564] <= 1'h0;
      write_done_data_log_force[2565] <= 1'h0;
      write_done_data_log_force[2566] <= 1'h0;
      write_done_data_log_force[2567] <= 1'h0;
      write_done_data_log_force[2568] <= 1'h0;
      write_done_data_log_force[2569] <= 1'h0;
      write_done_data_log_force[2570] <= 1'h0;
      write_done_data_log_force[2571] <= 1'h0;
      write_done_data_log_force[2572] <= 1'h0;
      write_done_data_log_force[2573] <= 1'h0;
      write_done_data_log_force[2574] <= 1'h0;
      write_done_data_log_force[2575] <= 1'h0;
      write_done_data_log_force[2576] <= 1'h0;
      write_done_data_log_force[2577] <= 1'h0;
      write_done_data_log_force[2578] <= 1'h0;
      write_done_data_log_force[2579] <= 1'h0;
      write_done_data_log_force[2580] <= 1'h0;
      write_done_data_log_force[2581] <= 1'h0;
      write_done_data_log_force[2582] <= 1'h0;
      write_done_data_log_force[2583] <= 1'h0;
      write_done_data_log_force[2584] <= 1'h0;
      write_done_data_log_force[2585] <= 1'h0;
      write_done_data_log_force[2586] <= 1'h0;
      write_done_data_log_force[2587] <= 1'h0;
      write_done_data_log_force[2588] <= 1'h0;
      write_done_data_log_force[2589] <= 1'h0;
      write_done_data_log_force[2590] <= 1'h0;
      write_done_data_log_force[2591] <= 1'h0;
      write_done_data_log_force[2592] <= 1'h0;
      write_done_data_log_force[2593] <= 1'h0;
      write_done_data_log_force[2594] <= 1'h0;
      write_done_data_log_force[2595] <= 1'h0;
      write_done_data_log_force[2596] <= 1'h0;
      write_done_data_log_force[2597] <= 1'h0;
      write_done_data_log_force[2598] <= 1'h0;
      write_done_data_log_force[2599] <= 1'h0;
      write_done_data_log_force[2600] <= 1'h0;
      write_done_data_log_force[2601] <= 1'h0;
      write_done_data_log_force[2602] <= 1'h0;
      write_done_data_log_force[2603] <= 1'h0;
      write_done_data_log_force[2604] <= 1'h0;
      write_done_data_log_force[2605] <= 1'h0;
      write_done_data_log_force[2606] <= 1'h0;
      write_done_data_log_force[2607] <= 1'h0;
      write_done_data_log_force[2608] <= 1'h0;
      write_done_data_log_force[2609] <= 1'h0;
      write_done_data_log_force[2610] <= 1'h0;
      write_done_data_log_force[2611] <= 1'h0;
      write_done_data_log_force[2612] <= 1'h0;
      write_done_data_log_force[2613] <= 1'h0;
      write_done_data_log_force[2614] <= 1'h0;
      write_done_data_log_force[2615] <= 1'h0;
      write_done_data_log_force[2616] <= 1'h0;
      write_done_data_log_force[2617] <= 1'h0;
      write_done_data_log_force[2618] <= 1'h0;
      write_done_data_log_force[2619] <= 1'h0;
      write_done_data_log_force[2620] <= 1'h0;
      write_done_data_log_force[2621] <= 1'h0;
      write_done_data_log_force[2622] <= 1'h0;
      write_done_data_log_force[2623] <= 1'h0;
      write_done_data_log_force[2624] <= 1'h0;
      write_done_data_log_force[2625] <= 1'h0;
      write_done_data_log_force[2626] <= 1'h0;
      write_done_data_log_force[2627] <= 1'h0;
      write_done_data_log_force[2628] <= 1'h0;
      write_done_data_log_force[2629] <= 1'h0;
      write_done_data_log_force[2630] <= 1'h0;
      write_done_data_log_force[2631] <= 1'h0;
      write_done_data_log_force[2632] <= 1'h0;
      write_done_data_log_force[2633] <= 1'h0;
      write_done_data_log_force[2634] <= 1'h0;
      write_done_data_log_force[2635] <= 1'h0;
      write_done_data_log_force[2636] <= 1'h0;
      write_done_data_log_force[2637] <= 1'h0;
      write_done_data_log_force[2638] <= 1'h0;
      write_done_data_log_force[2639] <= 1'h0;
      write_done_data_log_force[2640] <= 1'h0;
      write_done_data_log_force[2641] <= 1'h0;
      write_done_data_log_force[2642] <= 1'h0;
      write_done_data_log_force[2643] <= 1'h0;
      write_done_data_log_force[2644] <= 1'h0;
      write_done_data_log_force[2645] <= 1'h0;
      write_done_data_log_force[2646] <= 1'h0;
      write_done_data_log_force[2647] <= 1'h0;
      write_done_data_log_force[2648] <= 1'h0;
      write_done_data_log_force[2649] <= 1'h0;
      write_done_data_log_force[2650] <= 1'h0;
      write_done_data_log_force[2651] <= 1'h0;
      write_done_data_log_force[2652] <= 1'h0;
      write_done_data_log_force[2653] <= 1'h0;
      write_done_data_log_force[2654] <= 1'h0;
      write_done_data_log_force[2655] <= 1'h0;
      write_done_data_log_force[2656] <= 1'h0;
      write_done_data_log_force[2657] <= 1'h0;
      write_done_data_log_force[2658] <= 1'h0;
      write_done_data_log_force[2659] <= 1'h0;
      write_done_data_log_force[2660] <= 1'h0;
      write_done_data_log_force[2661] <= 1'h0;
      write_done_data_log_force[2662] <= 1'h0;
      write_done_data_log_force[2663] <= 1'h0;
      write_done_data_log_force[2664] <= 1'h0;
      write_done_data_log_force[2665] <= 1'h0;
      write_done_data_log_force[2666] <= 1'h0;
      write_done_data_log_force[2667] <= 1'h0;
      write_done_data_log_force[2668] <= 1'h0;
      write_done_data_log_force[2669] <= 1'h0;
      write_done_data_log_force[2670] <= 1'h0;
      write_done_data_log_force[2671] <= 1'h0;
      write_done_data_log_force[2672] <= 1'h0;
      write_done_data_log_force[2673] <= 1'h0;
      write_done_data_log_force[2674] <= 1'h0;
      write_done_data_log_force[2675] <= 1'h0;
      write_done_data_log_force[2676] <= 1'h0;
      write_done_data_log_force[2677] <= 1'h0;
      write_done_data_log_force[2678] <= 1'h0;
      write_done_data_log_force[2679] <= 1'h0;
      write_done_data_log_force[2680] <= 1'h0;
      write_done_data_log_force[2681] <= 1'h0;
      write_done_data_log_force[2682] <= 1'h0;
      write_done_data_log_force[2683] <= 1'h0;
      write_done_data_log_force[2684] <= 1'h0;
      write_done_data_log_force[2685] <= 1'h0;
      write_done_data_log_force[2686] <= 1'h0;
      write_done_data_log_force[2687] <= 1'h0;
      write_done_data_log_force[2688] <= 1'h0;
      write_done_data_log_force[2689] <= 1'h0;
      write_done_data_log_force[2690] <= 1'h0;
      write_done_data_log_force[2691] <= 1'h0;
      write_done_data_log_force[2692] <= 1'h0;
      write_done_data_log_force[2693] <= 1'h0;
      write_done_data_log_force[2694] <= 1'h0;
      write_done_data_log_force[2695] <= 1'h0;
      write_done_data_log_force[2696] <= 1'h0;
      write_done_data_log_force[2697] <= 1'h0;
      write_done_data_log_force[2698] <= 1'h0;
      write_done_data_log_force[2699] <= 1'h0;
      write_done_data_log_force[2700] <= 1'h0;
      write_done_data_log_force[2701] <= 1'h0;
      write_done_data_log_force[2702] <= 1'h0;
      write_done_data_log_force[2703] <= 1'h0;
      write_done_data_log_force[2704] <= 1'h0;
      write_done_data_log_force[2705] <= 1'h0;
      write_done_data_log_force[2706] <= 1'h0;
      write_done_data_log_force[2707] <= 1'h0;
      write_done_data_log_force[2708] <= 1'h0;
      write_done_data_log_force[2709] <= 1'h0;
      write_done_data_log_force[2710] <= 1'h0;
      write_done_data_log_force[2711] <= 1'h0;
      write_done_data_log_force[2712] <= 1'h0;
      write_done_data_log_force[2713] <= 1'h0;
      write_done_data_log_force[2714] <= 1'h0;
      write_done_data_log_force[2715] <= 1'h0;
      write_done_data_log_force[2716] <= 1'h0;
      write_done_data_log_force[2717] <= 1'h0;
      write_done_data_log_force[2718] <= 1'h0;
      write_done_data_log_force[2719] <= 1'h0;
      write_done_data_log_force[2720] <= 1'h0;
      write_done_data_log_force[2721] <= 1'h0;
      write_done_data_log_force[2722] <= 1'h0;
      write_done_data_log_force[2723] <= 1'h0;
      write_done_data_log_force[2724] <= 1'h0;
      write_done_data_log_force[2725] <= 1'h0;
      write_done_data_log_force[2726] <= 1'h0;
      write_done_data_log_force[2727] <= 1'h0;
      write_done_data_log_force[2728] <= 1'h0;
      write_done_data_log_force[2729] <= 1'h0;
      write_done_data_log_force[2730] <= 1'h0;
      write_done_data_log_force[2731] <= 1'h0;
      write_done_data_log_force[2732] <= 1'h0;
      write_done_data_log_force[2733] <= 1'h0;
      write_done_data_log_force[2734] <= 1'h0;
      write_done_data_log_force[2735] <= 1'h0;
      write_done_data_log_force[2736] <= 1'h0;
      write_done_data_log_force[2737] <= 1'h0;
      write_done_data_log_force[2738] <= 1'h0;
      write_done_data_log_force[2739] <= 1'h0;
      write_done_data_log_force[2740] <= 1'h0;
      write_done_data_log_force[2741] <= 1'h0;
      write_done_data_log_force[2742] <= 1'h0;
      write_done_data_log_force[2743] <= 1'h0;
      write_done_data_log_force[2744] <= 1'h0;
      write_done_data_log_force[2745] <= 1'h0;
      write_done_data_log_force[2746] <= 1'h0;
      write_done_data_log_force[2747] <= 1'h0;
      write_done_data_log_force[2748] <= 1'h0;
      write_done_data_log_force[2749] <= 1'h0;
      write_done_data_log_force[2750] <= 1'h0;
      write_done_data_log_force[2751] <= 1'h0;
      write_done_data_log_force[2752] <= 1'h0;
      write_done_data_log_force[2753] <= 1'h0;
      write_done_data_log_force[2754] <= 1'h0;
      write_done_data_log_force[2755] <= 1'h0;
      write_done_data_log_force[2756] <= 1'h0;
      write_done_data_log_force[2757] <= 1'h0;
      write_done_data_log_force[2758] <= 1'h0;
      write_done_data_log_force[2759] <= 1'h0;
      write_done_data_log_force[2760] <= 1'h0;
      write_done_data_log_force[2761] <= 1'h0;
      write_done_data_log_force[2762] <= 1'h0;
      write_done_data_log_force[2763] <= 1'h0;
      write_done_data_log_force[2764] <= 1'h0;
      write_done_data_log_force[2765] <= 1'h0;
      write_done_data_log_force[2766] <= 1'h0;
      write_done_data_log_force[2767] <= 1'h0;
      write_done_data_log_force[2768] <= 1'h0;
      write_done_data_log_force[2769] <= 1'h0;
      write_done_data_log_force[2770] <= 1'h0;
      write_done_data_log_force[2771] <= 1'h0;
      write_done_data_log_force[2772] <= 1'h0;
      write_done_data_log_force[2773] <= 1'h0;
      write_done_data_log_force[2774] <= 1'h0;
      write_done_data_log_force[2775] <= 1'h0;
      write_done_data_log_force[2776] <= 1'h0;
      write_done_data_log_force[2777] <= 1'h0;
      write_done_data_log_force[2778] <= 1'h0;
      write_done_data_log_force[2779] <= 1'h0;
      write_done_data_log_force[2780] <= 1'h0;
      write_done_data_log_force[2781] <= 1'h0;
      write_done_data_log_force[2782] <= 1'h0;
      write_done_data_log_force[2783] <= 1'h0;
      write_done_data_log_force[2784] <= 1'h0;
      write_done_data_log_force[2785] <= 1'h0;
      write_done_data_log_force[2786] <= 1'h0;
      write_done_data_log_force[2787] <= 1'h0;
      write_done_data_log_force[2788] <= 1'h0;
      write_done_data_log_force[2789] <= 1'h0;
      write_done_data_log_force[2790] <= 1'h0;
      write_done_data_log_force[2791] <= 1'h0;
      write_done_data_log_force[2792] <= 1'h0;
      write_done_data_log_force[2793] <= 1'h0;
      write_done_data_log_force[2794] <= 1'h0;
      write_done_data_log_force[2795] <= 1'h0;
      write_done_data_log_force[2796] <= 1'h0;
      write_done_data_log_force[2797] <= 1'h0;
      write_done_data_log_force[2798] <= 1'h0;
      write_done_data_log_force[2799] <= 1'h0;
      write_done_data_log_force[2800] <= 1'h0;
      write_done_data_log_force[2801] <= 1'h0;
      write_done_data_log_force[2802] <= 1'h0;
      write_done_data_log_force[2803] <= 1'h0;
      write_done_data_log_force[2804] <= 1'h0;
      write_done_data_log_force[2805] <= 1'h0;
      write_done_data_log_force[2806] <= 1'h0;
      write_done_data_log_force[2807] <= 1'h0;
      write_done_data_log_force[2808] <= 1'h0;
      write_done_data_log_force[2809] <= 1'h0;
      write_done_data_log_force[2810] <= 1'h0;
      write_done_data_log_force[2811] <= 1'h0;
      write_done_data_log_force[2812] <= 1'h0;
      write_done_data_log_force[2813] <= 1'h0;
      write_done_data_log_force[2814] <= 1'h0;
      write_done_data_log_force[2815] <= 1'h0;
      write_done_data_log_force[2816] <= 1'h0;
      write_done_data_log_force[2817] <= 1'h0;
      write_done_data_log_force[2818] <= 1'h0;
      write_done_data_log_force[2819] <= 1'h0;
      write_done_data_log_force[2820] <= 1'h0;
      write_done_data_log_force[2821] <= 1'h0;
      write_done_data_log_force[2822] <= 1'h0;
      write_done_data_log_force[2823] <= 1'h0;
      write_done_data_log_force[2824] <= 1'h0;
      write_done_data_log_force[2825] <= 1'h0;
      write_done_data_log_force[2826] <= 1'h0;
      write_done_data_log_force[2827] <= 1'h0;
      write_done_data_log_force[2828] <= 1'h0;
      write_done_data_log_force[2829] <= 1'h0;
      write_done_data_log_force[2830] <= 1'h0;
      write_done_data_log_force[2831] <= 1'h0;
      write_done_data_log_force[2832] <= 1'h0;
      write_done_data_log_force[2833] <= 1'h0;
      write_done_data_log_force[2834] <= 1'h0;
      write_done_data_log_force[2835] <= 1'h0;
      write_done_data_log_force[2836] <= 1'h0;
      write_done_data_log_force[2837] <= 1'h0;
      write_done_data_log_force[2838] <= 1'h0;
      write_done_data_log_force[2839] <= 1'h0;
      write_done_data_log_force[2840] <= 1'h0;
      write_done_data_log_force[2841] <= 1'h0;
      write_done_data_log_force[2842] <= 1'h0;
      write_done_data_log_force[2843] <= 1'h0;
      write_done_data_log_force[2844] <= 1'h0;
      write_done_data_log_force[2845] <= 1'h0;
      write_done_data_log_force[2846] <= 1'h0;
      write_done_data_log_force[2847] <= 1'h0;
      write_done_data_log_force[2848] <= 1'h0;
      write_done_data_log_force[2849] <= 1'h0;
      write_done_data_log_force[2850] <= 1'h0;
      write_done_data_log_force[2851] <= 1'h0;
      write_done_data_log_force[2852] <= 1'h0;
      write_done_data_log_force[2853] <= 1'h0;
      write_done_data_log_force[2854] <= 1'h0;
      write_done_data_log_force[2855] <= 1'h0;
      write_done_data_log_force[2856] <= 1'h0;
      write_done_data_log_force[2857] <= 1'h0;
      write_done_data_log_force[2858] <= 1'h0;
      write_done_data_log_force[2859] <= 1'h0;
      write_done_data_log_force[2860] <= 1'h0;
      write_done_data_log_force[2861] <= 1'h0;
      write_done_data_log_force[2862] <= 1'h0;
      write_done_data_log_force[2863] <= 1'h0;
      write_done_data_log_force[2864] <= 1'h0;
      write_done_data_log_force[2865] <= 1'h0;
      write_done_data_log_force[2866] <= 1'h0;
      write_done_data_log_force[2867] <= 1'h0;
      write_done_data_log_force[2868] <= 1'h0;
      write_done_data_log_force[2869] <= 1'h0;
      write_done_data_log_force[2870] <= 1'h0;
      write_done_data_log_force[2871] <= 1'h0;
      write_done_data_log_force[2872] <= 1'h0;
      write_done_data_log_force[2873] <= 1'h0;
      write_done_data_log_force[2874] <= 1'h0;
      write_done_data_log_force[2875] <= 1'h0;
      write_done_data_log_force[2876] <= 1'h0;
      write_done_data_log_force[2877] <= 1'h0;
      write_done_data_log_force[2878] <= 1'h0;
      write_done_data_log_force[2879] <= 1'h0;
      write_done_data_log_force[2880] <= 1'h0;
      write_done_data_log_force[2881] <= 1'h0;
      write_done_data_log_force[2882] <= 1'h0;
      write_done_data_log_force[2883] <= 1'h0;
      write_done_data_log_force[2884] <= 1'h0;
      write_done_data_log_force[2885] <= 1'h0;
      write_done_data_log_force[2886] <= 1'h0;
      write_done_data_log_force[2887] <= 1'h0;
      write_done_data_log_force[2888] <= 1'h0;
      write_done_data_log_force[2889] <= 1'h0;
      write_done_data_log_force[2890] <= 1'h0;
      write_done_data_log_force[2891] <= 1'h0;
      write_done_data_log_force[2892] <= 1'h0;
      write_done_data_log_force[2893] <= 1'h0;
      write_done_data_log_force[2894] <= 1'h0;
      write_done_data_log_force[2895] <= 1'h0;
      write_done_data_log_force[2896] <= 1'h0;
      write_done_data_log_force[2897] <= 1'h0;
      write_done_data_log_force[2898] <= 1'h0;
      write_done_data_log_force[2899] <= 1'h0;
      write_done_data_log_force[2900] <= 1'h0;
      write_done_data_log_force[2901] <= 1'h0;
      write_done_data_log_force[2902] <= 1'h0;
      write_done_data_log_force[2903] <= 1'h0;
      write_done_data_log_force[2904] <= 1'h0;
      write_done_data_log_force[2905] <= 1'h0;
      write_done_data_log_force[2906] <= 1'h0;
      write_done_data_log_force[2907] <= 1'h0;
      write_done_data_log_force[2908] <= 1'h0;
      write_done_data_log_force[2909] <= 1'h0;
      write_done_data_log_force[2910] <= 1'h0;
      write_done_data_log_force[2911] <= 1'h0;
      write_done_data_log_force[2912] <= 1'h0;
      write_done_data_log_force[2913] <= 1'h0;
      write_done_data_log_force[2914] <= 1'h0;
      write_done_data_log_force[2915] <= 1'h0;
      write_done_data_log_force[2916] <= 1'h0;
      write_done_data_log_force[2917] <= 1'h0;
      write_done_data_log_force[2918] <= 1'h0;
      write_done_data_log_force[2919] <= 1'h0;
      write_done_data_log_force[2920] <= 1'h0;
      write_done_data_log_force[2921] <= 1'h0;
      write_done_data_log_force[2922] <= 1'h0;
      write_done_data_log_force[2923] <= 1'h0;
      write_done_data_log_force[2924] <= 1'h0;
      write_done_data_log_force[2925] <= 1'h0;
      write_done_data_log_force[2926] <= 1'h0;
      write_done_data_log_force[2927] <= 1'h0;
      write_done_data_log_force[2928] <= 1'h0;
      write_done_data_log_force[2929] <= 1'h0;
      write_done_data_log_force[2930] <= 1'h0;
      write_done_data_log_force[2931] <= 1'h0;
      write_done_data_log_force[2932] <= 1'h0;
      write_done_data_log_force[2933] <= 1'h0;
      write_done_data_log_force[2934] <= 1'h0;
      write_done_data_log_force[2935] <= 1'h0;
      write_done_data_log_force[2936] <= 1'h0;
      write_done_data_log_force[2937] <= 1'h0;
      write_done_data_log_force[2938] <= 1'h0;
      write_done_data_log_force[2939] <= 1'h0;
      write_done_data_log_force[2940] <= 1'h0;
      write_done_data_log_force[2941] <= 1'h0;
      write_done_data_log_force[2942] <= 1'h0;
      write_done_data_log_force[2943] <= 1'h0;
      write_done_data_log_force[2944] <= 1'h0;
      write_done_data_log_force[2945] <= 1'h0;
      write_done_data_log_force[2946] <= 1'h0;
      write_done_data_log_force[2947] <= 1'h0;
      write_done_data_log_force[2948] <= 1'h0;
      write_done_data_log_force[2949] <= 1'h0;
      write_done_data_log_force[2950] <= 1'h0;
      write_done_data_log_force[2951] <= 1'h0;
      write_done_data_log_force[2952] <= 1'h0;
      write_done_data_log_force[2953] <= 1'h0;
      write_done_data_log_force[2954] <= 1'h0;
      write_done_data_log_force[2955] <= 1'h0;
      write_done_data_log_force[2956] <= 1'h0;
      write_done_data_log_force[2957] <= 1'h0;
      write_done_data_log_force[2958] <= 1'h0;
      write_done_data_log_force[2959] <= 1'h0;
      write_done_data_log_force[2960] <= 1'h0;
      write_done_data_log_force[2961] <= 1'h0;
      write_done_data_log_force[2962] <= 1'h0;
      write_done_data_log_force[2963] <= 1'h0;
      write_done_data_log_force[2964] <= 1'h0;
      write_done_data_log_force[2965] <= 1'h0;
      write_done_data_log_force[2966] <= 1'h0;
      write_done_data_log_force[2967] <= 1'h0;
      write_done_data_log_force[2968] <= 1'h0;
      write_done_data_log_force[2969] <= 1'h0;
      write_done_data_log_force[2970] <= 1'h0;
      write_done_data_log_force[2971] <= 1'h0;
      write_done_data_log_force[2972] <= 1'h0;
      write_done_data_log_force[2973] <= 1'h0;
      write_done_data_log_force[2974] <= 1'h0;
      write_done_data_log_force[2975] <= 1'h0;
      write_done_data_log_force[2976] <= 1'h0;
      write_done_data_log_force[2977] <= 1'h0;
      write_done_data_log_force[2978] <= 1'h0;
      write_done_data_log_force[2979] <= 1'h0;
      write_done_data_log_force[2980] <= 1'h0;
      write_done_data_log_force[2981] <= 1'h0;
      write_done_data_log_force[2982] <= 1'h0;
      write_done_data_log_force[2983] <= 1'h0;
      write_done_data_log_force[2984] <= 1'h0;
      write_done_data_log_force[2985] <= 1'h0;
      write_done_data_log_force[2986] <= 1'h0;
      write_done_data_log_force[2987] <= 1'h0;
      write_done_data_log_force[2988] <= 1'h0;
      write_done_data_log_force[2989] <= 1'h0;
      write_done_data_log_force[2990] <= 1'h0;
      write_done_data_log_force[2991] <= 1'h0;
      write_done_data_log_force[2992] <= 1'h0;
      write_done_data_log_force[2993] <= 1'h0;
      write_done_data_log_force[2994] <= 1'h0;
      write_done_data_log_force[2995] <= 1'h0;
      write_done_data_log_force[2996] <= 1'h0;
      write_done_data_log_force[2997] <= 1'h0;
      write_done_data_log_force[2998] <= 1'h0;
      write_done_data_log_force[2999] <= 1'h0;
      write_done_data_log_force[3000] <= 1'h0;
      write_done_data_log_force[3001] <= 1'h0;
      write_done_data_log_force[3002] <= 1'h0;
      write_done_data_log_force[3003] <= 1'h0;
      write_done_data_log_force[3004] <= 1'h0;
      write_done_data_log_force[3005] <= 1'h0;
      write_done_data_log_force[3006] <= 1'h0;
      write_done_data_log_force[3007] <= 1'h0;
      write_done_data_log_force[3008] <= 1'h0;
      write_done_data_log_force[3009] <= 1'h0;
      write_done_data_log_force[3010] <= 1'h0;
      write_done_data_log_force[3011] <= 1'h0;
      write_done_data_log_force[3012] <= 1'h0;
      write_done_data_log_force[3013] <= 1'h0;
      write_done_data_log_force[3014] <= 1'h0;
      write_done_data_log_force[3015] <= 1'h0;
      write_done_data_log_force[3016] <= 1'h0;
      write_done_data_log_force[3017] <= 1'h0;
      write_done_data_log_force[3018] <= 1'h0;
      write_done_data_log_force[3019] <= 1'h0;
      write_done_data_log_force[3020] <= 1'h0;
      write_done_data_log_force[3021] <= 1'h0;
      write_done_data_log_force[3022] <= 1'h0;
      write_done_data_log_force[3023] <= 1'h0;
      write_done_data_log_force[3024] <= 1'h0;
      write_done_data_log_force[3025] <= 1'h0;
      write_done_data_log_force[3026] <= 1'h0;
      write_done_data_log_force[3027] <= 1'h0;
      write_done_data_log_force[3028] <= 1'h0;
      write_done_data_log_force[3029] <= 1'h0;
      write_done_data_log_force[3030] <= 1'h0;
      write_done_data_log_force[3031] <= 1'h0;
      write_done_data_log_force[3032] <= 1'h0;
      write_done_data_log_force[3033] <= 1'h0;
      write_done_data_log_force[3034] <= 1'h0;
      write_done_data_log_force[3035] <= 1'h0;
      write_done_data_log_force[3036] <= 1'h0;
      write_done_data_log_force[3037] <= 1'h0;
      write_done_data_log_force[3038] <= 1'h0;
      write_done_data_log_force[3039] <= 1'h0;
      write_done_data_log_force[3040] <= 1'h0;
      write_done_data_log_force[3041] <= 1'h0;
      write_done_data_log_force[3042] <= 1'h0;
      write_done_data_log_force[3043] <= 1'h0;
      write_done_data_log_force[3044] <= 1'h0;
      write_done_data_log_force[3045] <= 1'h0;
      write_done_data_log_force[3046] <= 1'h0;
      write_done_data_log_force[3047] <= 1'h0;
      write_done_data_log_force[3048] <= 1'h0;
      write_done_data_log_force[3049] <= 1'h0;
      write_done_data_log_force[3050] <= 1'h0;
      write_done_data_log_force[3051] <= 1'h0;
      write_done_data_log_force[3052] <= 1'h0;
      write_done_data_log_force[3053] <= 1'h0;
      write_done_data_log_force[3054] <= 1'h0;
      write_done_data_log_force[3055] <= 1'h0;
      write_done_data_log_force[3056] <= 1'h0;
      write_done_data_log_force[3057] <= 1'h0;
      write_done_data_log_force[3058] <= 1'h0;
      write_done_data_log_force[3059] <= 1'h0;
      write_done_data_log_force[3060] <= 1'h0;
      write_done_data_log_force[3061] <= 1'h0;
      write_done_data_log_force[3062] <= 1'h0;
      write_done_data_log_force[3063] <= 1'h0;
      write_done_data_log_force[3064] <= 1'h0;
      write_done_data_log_force[3065] <= 1'h0;
      write_done_data_log_force[3066] <= 1'h0;
      write_done_data_log_force[3067] <= 1'h0;
      write_done_data_log_force[3068] <= 1'h0;
      write_done_data_log_force[3069] <= 1'h0;
      write_done_data_log_force[3070] <= 1'h0;
      write_done_data_log_force[3071] <= 1'h0;
      write_done_data_log_force[3072] <= 1'h0;
      write_done_data_log_force[3073] <= 1'h0;
      write_done_data_log_force[3074] <= 1'h0;
      write_done_data_log_force[3075] <= 1'h0;
      write_done_data_log_force[3076] <= 1'h0;
      write_done_data_log_force[3077] <= 1'h0;
      write_done_data_log_force[3078] <= 1'h0;
      write_done_data_log_force[3079] <= 1'h0;
      write_done_data_log_force[3080] <= 1'h0;
      write_done_data_log_force[3081] <= 1'h0;
      write_done_data_log_force[3082] <= 1'h0;
      write_done_data_log_force[3083] <= 1'h0;
      write_done_data_log_force[3084] <= 1'h0;
      write_done_data_log_force[3085] <= 1'h0;
      write_done_data_log_force[3086] <= 1'h0;
      write_done_data_log_force[3087] <= 1'h0;
      write_done_data_log_force[3088] <= 1'h0;
      write_done_data_log_force[3089] <= 1'h0;
      write_done_data_log_force[3090] <= 1'h0;
      write_done_data_log_force[3091] <= 1'h0;
      write_done_data_log_force[3092] <= 1'h0;
      write_done_data_log_force[3093] <= 1'h0;
      write_done_data_log_force[3094] <= 1'h0;
      write_done_data_log_force[3095] <= 1'h0;
      write_done_data_log_force[3096] <= 1'h0;
      write_done_data_log_force[3097] <= 1'h0;
      write_done_data_log_force[3098] <= 1'h0;
      write_done_data_log_force[3099] <= 1'h0;
      write_done_data_log_force[3100] <= 1'h0;
      write_done_data_log_force[3101] <= 1'h0;
      write_done_data_log_force[3102] <= 1'h0;
      write_done_data_log_force[3103] <= 1'h0;
      write_done_data_log_force[3104] <= 1'h0;
      write_done_data_log_force[3105] <= 1'h0;
      write_done_data_log_force[3106] <= 1'h0;
      write_done_data_log_force[3107] <= 1'h0;
      write_done_data_log_force[3108] <= 1'h0;
      write_done_data_log_force[3109] <= 1'h0;
      write_done_data_log_force[3110] <= 1'h0;
      write_done_data_log_force[3111] <= 1'h0;
      write_done_data_log_force[3112] <= 1'h0;
      write_done_data_log_force[3113] <= 1'h0;
      write_done_data_log_force[3114] <= 1'h0;
      write_done_data_log_force[3115] <= 1'h0;
      write_done_data_log_force[3116] <= 1'h0;
      write_done_data_log_force[3117] <= 1'h0;
      write_done_data_log_force[3118] <= 1'h0;
      write_done_data_log_force[3119] <= 1'h0;
      write_done_data_log_force[3120] <= 1'h0;
      write_done_data_log_force[3121] <= 1'h0;
      write_done_data_log_force[3122] <= 1'h0;
      write_done_data_log_force[3123] <= 1'h0;
      write_done_data_log_force[3124] <= 1'h0;
      write_done_data_log_force[3125] <= 1'h0;
      write_done_data_log_force[3126] <= 1'h0;
      write_done_data_log_force[3127] <= 1'h0;
      write_done_data_log_force[3128] <= 1'h0;
      write_done_data_log_force[3129] <= 1'h0;
      write_done_data_log_force[3130] <= 1'h0;
      write_done_data_log_force[3131] <= 1'h0;
      write_done_data_log_force[3132] <= 1'h0;
      write_done_data_log_force[3133] <= 1'h0;
      write_done_data_log_force[3134] <= 1'h0;
      write_done_data_log_force[3135] <= 1'h0;
      write_done_data_log_force[3136] <= 1'h0;
      write_done_data_log_force[3137] <= 1'h0;
      write_done_data_log_force[3138] <= 1'h0;
      write_done_data_log_force[3139] <= 1'h0;
      write_done_data_log_force[3140] <= 1'h0;
      write_done_data_log_force[3141] <= 1'h0;
      write_done_data_log_force[3142] <= 1'h0;
      write_done_data_log_force[3143] <= 1'h0;
      write_done_data_log_force[3144] <= 1'h0;
      write_done_data_log_force[3145] <= 1'h0;
      write_done_data_log_force[3146] <= 1'h0;
      write_done_data_log_force[3147] <= 1'h0;
      write_done_data_log_force[3148] <= 1'h0;
      write_done_data_log_force[3149] <= 1'h0;
      write_done_data_log_force[3150] <= 1'h0;
      write_done_data_log_force[3151] <= 1'h0;
      write_done_data_log_force[3152] <= 1'h0;
      write_done_data_log_force[3153] <= 1'h0;
      write_done_data_log_force[3154] <= 1'h0;
      write_done_data_log_force[3155] <= 1'h0;
      write_done_data_log_force[3156] <= 1'h0;
      write_done_data_log_force[3157] <= 1'h0;
      write_done_data_log_force[3158] <= 1'h0;
      write_done_data_log_force[3159] <= 1'h0;
      write_done_data_log_force[3160] <= 1'h0;
      write_done_data_log_force[3161] <= 1'h0;
      write_done_data_log_force[3162] <= 1'h0;
      write_done_data_log_force[3163] <= 1'h0;
      write_done_data_log_force[3164] <= 1'h0;
      write_done_data_log_force[3165] <= 1'h0;
      write_done_data_log_force[3166] <= 1'h0;
      write_done_data_log_force[3167] <= 1'h0;
      write_done_data_log_force[3168] <= 1'h0;
      write_done_data_log_force[3169] <= 1'h0;
      write_done_data_log_force[3170] <= 1'h0;
      write_done_data_log_force[3171] <= 1'h0;
      write_done_data_log_force[3172] <= 1'h0;
      write_done_data_log_force[3173] <= 1'h0;
      write_done_data_log_force[3174] <= 1'h0;
      write_done_data_log_force[3175] <= 1'h0;
      write_done_data_log_force[3176] <= 1'h0;
      write_done_data_log_force[3177] <= 1'h0;
      write_done_data_log_force[3178] <= 1'h0;
      write_done_data_log_force[3179] <= 1'h0;
      write_done_data_log_force[3180] <= 1'h0;
      write_done_data_log_force[3181] <= 1'h0;
      write_done_data_log_force[3182] <= 1'h0;
      write_done_data_log_force[3183] <= 1'h0;
      write_done_data_log_force[3184] <= 1'h0;
      write_done_data_log_force[3185] <= 1'h0;
      write_done_data_log_force[3186] <= 1'h0;
      write_done_data_log_force[3187] <= 1'h0;
      write_done_data_log_force[3188] <= 1'h0;
      write_done_data_log_force[3189] <= 1'h0;
      write_done_data_log_force[3190] <= 1'h0;
      write_done_data_log_force[3191] <= 1'h0;
      write_done_data_log_force[3192] <= 1'h0;
      write_done_data_log_force[3193] <= 1'h0;
      write_done_data_log_force[3194] <= 1'h0;
      write_done_data_log_force[3195] <= 1'h0;
      write_done_data_log_force[3196] <= 1'h0;
      write_done_data_log_force[3197] <= 1'h0;
      write_done_data_log_force[3198] <= 1'h0;
      write_done_data_log_force[3199] <= 1'h0;
      write_done_data_log_force[3200] <= 1'h0;
      write_done_data_log_force[3201] <= 1'h0;
      write_done_data_log_force[3202] <= 1'h0;
      write_done_data_log_force[3203] <= 1'h0;
      write_done_data_log_force[3204] <= 1'h0;
      write_done_data_log_force[3205] <= 1'h0;
      write_done_data_log_force[3206] <= 1'h0;
      write_done_data_log_force[3207] <= 1'h0;
      write_done_data_log_force[3208] <= 1'h0;
      write_done_data_log_force[3209] <= 1'h0;
      write_done_data_log_force[3210] <= 1'h0;
      write_done_data_log_force[3211] <= 1'h0;
      write_done_data_log_force[3212] <= 1'h0;
      write_done_data_log_force[3213] <= 1'h0;
      write_done_data_log_force[3214] <= 1'h0;
      write_done_data_log_force[3215] <= 1'h0;
      write_done_data_log_force[3216] <= 1'h0;
      write_done_data_log_force[3217] <= 1'h0;
      write_done_data_log_force[3218] <= 1'h0;
      write_done_data_log_force[3219] <= 1'h0;
      write_done_data_log_force[3220] <= 1'h0;
      write_done_data_log_force[3221] <= 1'h0;
      write_done_data_log_force[3222] <= 1'h0;
      write_done_data_log_force[3223] <= 1'h0;
      write_done_data_log_force[3224] <= 1'h0;
      write_done_data_log_force[3225] <= 1'h0;
      write_done_data_log_force[3226] <= 1'h0;
      write_done_data_log_force[3227] <= 1'h0;
      write_done_data_log_force[3228] <= 1'h0;
      write_done_data_log_force[3229] <= 1'h0;
      write_done_data_log_force[3230] <= 1'h0;
      write_done_data_log_force[3231] <= 1'h0;
      write_done_data_log_force[3232] <= 1'h0;
      write_done_data_log_force[3233] <= 1'h0;
      write_done_data_log_force[3234] <= 1'h0;
      write_done_data_log_force[3235] <= 1'h0;
      write_done_data_log_force[3236] <= 1'h0;
      write_done_data_log_force[3237] <= 1'h0;
      write_done_data_log_force[3238] <= 1'h0;
      write_done_data_log_force[3239] <= 1'h0;
      write_done_data_log_force[3240] <= 1'h0;
      write_done_data_log_force[3241] <= 1'h0;
      write_done_data_log_force[3242] <= 1'h0;
      write_done_data_log_force[3243] <= 1'h0;
      write_done_data_log_force[3244] <= 1'h0;
      write_done_data_log_force[3245] <= 1'h0;
      write_done_data_log_force[3246] <= 1'h0;
      write_done_data_log_force[3247] <= 1'h0;
      write_done_data_log_force[3248] <= 1'h0;
      write_done_data_log_force[3249] <= 1'h0;
      write_done_data_log_force[3250] <= 1'h0;
      write_done_data_log_force[3251] <= 1'h0;
      write_done_data_log_force[3252] <= 1'h0;
      write_done_data_log_force[3253] <= 1'h0;
      write_done_data_log_force[3254] <= 1'h0;
      write_done_data_log_force[3255] <= 1'h0;
      write_done_data_log_force[3256] <= 1'h0;
      write_done_data_log_force[3257] <= 1'h0;
      write_done_data_log_force[3258] <= 1'h0;
      write_done_data_log_force[3259] <= 1'h0;
      write_done_data_log_force[3260] <= 1'h0;
      write_done_data_log_force[3261] <= 1'h0;
      write_done_data_log_force[3262] <= 1'h0;
      write_done_data_log_force[3263] <= 1'h0;
      write_done_data_log_force[3264] <= 1'h0;
      write_done_data_log_force[3265] <= 1'h0;
      write_done_data_log_force[3266] <= 1'h0;
      write_done_data_log_force[3267] <= 1'h0;
      write_done_data_log_force[3268] <= 1'h0;
      write_done_data_log_force[3269] <= 1'h0;
      write_done_data_log_force[3270] <= 1'h0;
      write_done_data_log_force[3271] <= 1'h0;
      write_done_data_log_force[3272] <= 1'h0;
      write_done_data_log_force[3273] <= 1'h0;
      write_done_data_log_force[3274] <= 1'h0;
      write_done_data_log_force[3275] <= 1'h0;
      write_done_data_log_force[3276] <= 1'h0;
      write_done_data_log_force[3277] <= 1'h0;
      write_done_data_log_force[3278] <= 1'h0;
      write_done_data_log_force[3279] <= 1'h0;
      write_done_data_log_force[3280] <= 1'h0;
      write_done_data_log_force[3281] <= 1'h0;
      write_done_data_log_force[3282] <= 1'h0;
      write_done_data_log_force[3283] <= 1'h0;
      write_done_data_log_force[3284] <= 1'h0;
      write_done_data_log_force[3285] <= 1'h0;
      write_done_data_log_force[3286] <= 1'h0;
      write_done_data_log_force[3287] <= 1'h0;
      write_done_data_log_force[3288] <= 1'h0;
      write_done_data_log_force[3289] <= 1'h0;
      write_done_data_log_force[3290] <= 1'h0;
      write_done_data_log_force[3291] <= 1'h0;
      write_done_data_log_force[3292] <= 1'h0;
      write_done_data_log_force[3293] <= 1'h0;
      write_done_data_log_force[3294] <= 1'h0;
      write_done_data_log_force[3295] <= 1'h0;
      write_done_data_log_force[3296] <= 1'h0;
      write_done_data_log_force[3297] <= 1'h0;
      write_done_data_log_force[3298] <= 1'h0;
      write_done_data_log_force[3299] <= 1'h0;
      write_done_data_log_force[3300] <= 1'h0;
      write_done_data_log_force[3301] <= 1'h0;
      write_done_data_log_force[3302] <= 1'h0;
      write_done_data_log_force[3303] <= 1'h0;
      write_done_data_log_force[3304] <= 1'h0;
      write_done_data_log_force[3305] <= 1'h0;
      write_done_data_log_force[3306] <= 1'h0;
      write_done_data_log_force[3307] <= 1'h0;
      write_done_data_log_force[3308] <= 1'h0;
      write_done_data_log_force[3309] <= 1'h0;
      write_done_data_log_force[3310] <= 1'h0;
      write_done_data_log_force[3311] <= 1'h0;
      write_done_data_log_force[3312] <= 1'h0;
      write_done_data_log_force[3313] <= 1'h0;
      write_done_data_log_force[3314] <= 1'h0;
      write_done_data_log_force[3315] <= 1'h0;
      write_done_data_log_force[3316] <= 1'h0;
      write_done_data_log_force[3317] <= 1'h0;
      write_done_data_log_force[3318] <= 1'h0;
      write_done_data_log_force[3319] <= 1'h0;
      write_done_data_log_force[3320] <= 1'h0;
      write_done_data_log_force[3321] <= 1'h0;
      write_done_data_log_force[3322] <= 1'h0;
      write_done_data_log_force[3323] <= 1'h0;
      write_done_data_log_force[3324] <= 1'h0;
      write_done_data_log_force[3325] <= 1'h0;
      write_done_data_log_force[3326] <= 1'h0;
      write_done_data_log_force[3327] <= 1'h0;
      write_done_data_log_force[3328] <= 1'h0;
      write_done_data_log_force[3329] <= 1'h0;
      write_done_data_log_force[3330] <= 1'h0;
      write_done_data_log_force[3331] <= 1'h0;
      write_done_data_log_force[3332] <= 1'h0;
      write_done_data_log_force[3333] <= 1'h0;
      write_done_data_log_force[3334] <= 1'h0;
      write_done_data_log_force[3335] <= 1'h0;
      write_done_data_log_force[3336] <= 1'h0;
      write_done_data_log_force[3337] <= 1'h0;
      write_done_data_log_force[3338] <= 1'h0;
      write_done_data_log_force[3339] <= 1'h0;
      write_done_data_log_force[3340] <= 1'h0;
      write_done_data_log_force[3341] <= 1'h0;
      write_done_data_log_force[3342] <= 1'h0;
      write_done_data_log_force[3343] <= 1'h0;
      write_done_data_log_force[3344] <= 1'h0;
      write_done_data_log_force[3345] <= 1'h0;
      write_done_data_log_force[3346] <= 1'h0;
      write_done_data_log_force[3347] <= 1'h0;
      write_done_data_log_force[3348] <= 1'h0;
      write_done_data_log_force[3349] <= 1'h0;
      write_done_data_log_force[3350] <= 1'h0;
      write_done_data_log_force[3351] <= 1'h0;
      write_done_data_log_force[3352] <= 1'h0;
      write_done_data_log_force[3353] <= 1'h0;
      write_done_data_log_force[3354] <= 1'h0;
      write_done_data_log_force[3355] <= 1'h0;
      write_done_data_log_force[3356] <= 1'h0;
      write_done_data_log_force[3357] <= 1'h0;
      write_done_data_log_force[3358] <= 1'h0;
      write_done_data_log_force[3359] <= 1'h0;
      write_done_data_log_force[3360] <= 1'h0;
      write_done_data_log_force[3361] <= 1'h0;
      write_done_data_log_force[3362] <= 1'h0;
      write_done_data_log_force[3363] <= 1'h0;
      write_done_data_log_force[3364] <= 1'h0;
      write_done_data_log_force[3365] <= 1'h0;
      write_done_data_log_force[3366] <= 1'h0;
      write_done_data_log_force[3367] <= 1'h0;
      write_done_data_log_force[3368] <= 1'h0;
      write_done_data_log_force[3369] <= 1'h0;
      write_done_data_log_force[3370] <= 1'h0;
      write_done_data_log_force[3371] <= 1'h0;
      write_done_data_log_force[3372] <= 1'h0;
      write_done_data_log_force[3373] <= 1'h0;
      write_done_data_log_force[3374] <= 1'h0;
      write_done_data_log_force[3375] <= 1'h0;
      write_done_data_log_force[3376] <= 1'h0;
      write_done_data_log_force[3377] <= 1'h0;
      write_done_data_log_force[3378] <= 1'h0;
      write_done_data_log_force[3379] <= 1'h0;
      write_done_data_log_force[3380] <= 1'h0;
      write_done_data_log_force[3381] <= 1'h0;
      write_done_data_log_force[3382] <= 1'h0;
      write_done_data_log_force[3383] <= 1'h0;
      write_done_data_log_force[3384] <= 1'h0;
      write_done_data_log_force[3385] <= 1'h0;
      write_done_data_log_force[3386] <= 1'h0;
      write_done_data_log_force[3387] <= 1'h0;
      write_done_data_log_force[3388] <= 1'h0;
      write_done_data_log_force[3389] <= 1'h0;
      write_done_data_log_force[3390] <= 1'h0;
      write_done_data_log_force[3391] <= 1'h0;
      write_done_data_log_force[3392] <= 1'h0;
      write_done_data_log_force[3393] <= 1'h0;
      write_done_data_log_force[3394] <= 1'h0;
      write_done_data_log_force[3395] <= 1'h0;
      write_done_data_log_force[3396] <= 1'h0;
      write_done_data_log_force[3397] <= 1'h0;
      write_done_data_log_force[3398] <= 1'h0;
      write_done_data_log_force[3399] <= 1'h0;
      write_done_data_log_force[3400] <= 1'h0;
      write_done_data_log_force[3401] <= 1'h0;
      write_done_data_log_force[3402] <= 1'h0;
      write_done_data_log_force[3403] <= 1'h0;
      write_done_data_log_force[3404] <= 1'h0;
      write_done_data_log_force[3405] <= 1'h0;
      write_done_data_log_force[3406] <= 1'h0;
      write_done_data_log_force[3407] <= 1'h0;
      write_done_data_log_force[3408] <= 1'h0;
      write_done_data_log_force[3409] <= 1'h0;
      write_done_data_log_force[3410] <= 1'h0;
      write_done_data_log_force[3411] <= 1'h0;
      write_done_data_log_force[3412] <= 1'h0;
      write_done_data_log_force[3413] <= 1'h0;
      write_done_data_log_force[3414] <= 1'h0;
      write_done_data_log_force[3415] <= 1'h0;
      write_done_data_log_force[3416] <= 1'h0;
      write_done_data_log_force[3417] <= 1'h0;
      write_done_data_log_force[3418] <= 1'h0;
      write_done_data_log_force[3419] <= 1'h0;
      write_done_data_log_force[3420] <= 1'h0;
      write_done_data_log_force[3421] <= 1'h0;
      write_done_data_log_force[3422] <= 1'h0;
      write_done_data_log_force[3423] <= 1'h0;
      write_done_data_log_force[3424] <= 1'h0;
      write_done_data_log_force[3425] <= 1'h0;
      write_done_data_log_force[3426] <= 1'h0;
      write_done_data_log_force[3427] <= 1'h0;
      write_done_data_log_force[3428] <= 1'h0;
      write_done_data_log_force[3429] <= 1'h0;
      write_done_data_log_force[3430] <= 1'h0;
      write_done_data_log_force[3431] <= 1'h0;
      write_done_data_log_force[3432] <= 1'h0;
      write_done_data_log_force[3433] <= 1'h0;
      write_done_data_log_force[3434] <= 1'h0;
      write_done_data_log_force[3435] <= 1'h0;
      write_done_data_log_force[3436] <= 1'h0;
      write_done_data_log_force[3437] <= 1'h0;
      write_done_data_log_force[3438] <= 1'h0;
      write_done_data_log_force[3439] <= 1'h0;
      write_done_data_log_force[3440] <= 1'h0;
      write_done_data_log_force[3441] <= 1'h0;
      write_done_data_log_force[3442] <= 1'h0;
      write_done_data_log_force[3443] <= 1'h0;
      write_done_data_log_force[3444] <= 1'h0;
      write_done_data_log_force[3445] <= 1'h0;
      write_done_data_log_force[3446] <= 1'h0;
      write_done_data_log_force[3447] <= 1'h0;
      write_done_data_log_force[3448] <= 1'h0;
      write_done_data_log_force[3449] <= 1'h0;
      write_done_data_log_force[3450] <= 1'h0;
      write_done_data_log_force[3451] <= 1'h0;
      write_done_data_log_force[3452] <= 1'h0;
      write_done_data_log_force[3453] <= 1'h0;
      write_done_data_log_force[3454] <= 1'h0;
      write_done_data_log_force[3455] <= 1'h0;
      write_done_data_log_force[3456] <= 1'h0;
      write_done_data_log_force[3457] <= 1'h0;
      write_done_data_log_force[3458] <= 1'h0;
      write_done_data_log_force[3459] <= 1'h0;
      write_done_data_log_force[3460] <= 1'h0;
      write_done_data_log_force[3461] <= 1'h0;
      write_done_data_log_force[3462] <= 1'h0;
      write_done_data_log_force[3463] <= 1'h0;
      write_done_data_log_force[3464] <= 1'h0;
      write_done_data_log_force[3465] <= 1'h0;
      write_done_data_log_force[3466] <= 1'h0;
      write_done_data_log_force[3467] <= 1'h0;
      write_done_data_log_force[3468] <= 1'h0;
      write_done_data_log_force[3469] <= 1'h0;
      write_done_data_log_force[3470] <= 1'h0;
      write_done_data_log_force[3471] <= 1'h0;
      write_done_data_log_force[3472] <= 1'h0;
      write_done_data_log_force[3473] <= 1'h0;
      write_done_data_log_force[3474] <= 1'h0;
      write_done_data_log_force[3475] <= 1'h0;
      write_done_data_log_force[3476] <= 1'h0;
      write_done_data_log_force[3477] <= 1'h0;
      write_done_data_log_force[3478] <= 1'h0;
      write_done_data_log_force[3479] <= 1'h0;
      write_done_data_log_force[3480] <= 1'h0;
      write_done_data_log_force[3481] <= 1'h0;
      write_done_data_log_force[3482] <= 1'h0;
      write_done_data_log_force[3483] <= 1'h0;
      write_done_data_log_force[3484] <= 1'h0;
      write_done_data_log_force[3485] <= 1'h0;
      write_done_data_log_force[3486] <= 1'h0;
      write_done_data_log_force[3487] <= 1'h0;
      write_done_data_log_force[3488] <= 1'h0;
      write_done_data_log_force[3489] <= 1'h0;
      write_done_data_log_force[3490] <= 1'h0;
      write_done_data_log_force[3491] <= 1'h0;
      write_done_data_log_force[3492] <= 1'h0;
      write_done_data_log_force[3493] <= 1'h0;
      write_done_data_log_force[3494] <= 1'h0;
      write_done_data_log_force[3495] <= 1'h0;
      write_done_data_log_force[3496] <= 1'h0;
      write_done_data_log_force[3497] <= 1'h0;
      write_done_data_log_force[3498] <= 1'h0;
      write_done_data_log_force[3499] <= 1'h0;
      write_done_data_log_force[3500] <= 1'h0;
      write_done_data_log_force[3501] <= 1'h0;
      write_done_data_log_force[3502] <= 1'h0;
      write_done_data_log_force[3503] <= 1'h0;
      write_done_data_log_force[3504] <= 1'h0;
      write_done_data_log_force[3505] <= 1'h0;
      write_done_data_log_force[3506] <= 1'h0;
      write_done_data_log_force[3507] <= 1'h0;
      write_done_data_log_force[3508] <= 1'h0;
      write_done_data_log_force[3509] <= 1'h0;
      write_done_data_log_force[3510] <= 1'h0;
      write_done_data_log_force[3511] <= 1'h0;
      write_done_data_log_force[3512] <= 1'h0;
      write_done_data_log_force[3513] <= 1'h0;
      write_done_data_log_force[3514] <= 1'h0;
      write_done_data_log_force[3515] <= 1'h0;
      write_done_data_log_force[3516] <= 1'h0;
      write_done_data_log_force[3517] <= 1'h0;
      write_done_data_log_force[3518] <= 1'h0;
      write_done_data_log_force[3519] <= 1'h0;
      write_done_data_log_force[3520] <= 1'h0;
      write_done_data_log_force[3521] <= 1'h0;
      write_done_data_log_force[3522] <= 1'h0;
      write_done_data_log_force[3523] <= 1'h0;
      write_done_data_log_force[3524] <= 1'h0;
      write_done_data_log_force[3525] <= 1'h0;
      write_done_data_log_force[3526] <= 1'h0;
      write_done_data_log_force[3527] <= 1'h0;
      write_done_data_log_force[3528] <= 1'h0;
      write_done_data_log_force[3529] <= 1'h0;
      write_done_data_log_force[3530] <= 1'h0;
      write_done_data_log_force[3531] <= 1'h0;
      write_done_data_log_force[3532] <= 1'h0;
      write_done_data_log_force[3533] <= 1'h0;
      write_done_data_log_force[3534] <= 1'h0;
      write_done_data_log_force[3535] <= 1'h0;
      write_done_data_log_force[3536] <= 1'h0;
      write_done_data_log_force[3537] <= 1'h0;
      write_done_data_log_force[3538] <= 1'h0;
      write_done_data_log_force[3539] <= 1'h0;
      write_done_data_log_force[3540] <= 1'h0;
      write_done_data_log_force[3541] <= 1'h0;
      write_done_data_log_force[3542] <= 1'h0;
      write_done_data_log_force[3543] <= 1'h0;
      write_done_data_log_force[3544] <= 1'h0;
      write_done_data_log_force[3545] <= 1'h0;
      write_done_data_log_force[3546] <= 1'h0;
      write_done_data_log_force[3547] <= 1'h0;
      write_done_data_log_force[3548] <= 1'h0;
      write_done_data_log_force[3549] <= 1'h0;
      write_done_data_log_force[3550] <= 1'h0;
      write_done_data_log_force[3551] <= 1'h0;
      write_done_data_log_force[3552] <= 1'h0;
      write_done_data_log_force[3553] <= 1'h0;
      write_done_data_log_force[3554] <= 1'h0;
      write_done_data_log_force[3555] <= 1'h0;
      write_done_data_log_force[3556] <= 1'h0;
      write_done_data_log_force[3557] <= 1'h0;
      write_done_data_log_force[3558] <= 1'h0;
      write_done_data_log_force[3559] <= 1'h0;
      write_done_data_log_force[3560] <= 1'h0;
      write_done_data_log_force[3561] <= 1'h0;
      write_done_data_log_force[3562] <= 1'h0;
      write_done_data_log_force[3563] <= 1'h0;
      write_done_data_log_force[3564] <= 1'h0;
      write_done_data_log_force[3565] <= 1'h0;
      write_done_data_log_force[3566] <= 1'h0;
      write_done_data_log_force[3567] <= 1'h0;
      write_done_data_log_force[3568] <= 1'h0;
      write_done_data_log_force[3569] <= 1'h0;
      write_done_data_log_force[3570] <= 1'h0;
      write_done_data_log_force[3571] <= 1'h0;
      write_done_data_log_force[3572] <= 1'h0;
      write_done_data_log_force[3573] <= 1'h0;
      write_done_data_log_force[3574] <= 1'h0;
      write_done_data_log_force[3575] <= 1'h0;
      write_done_data_log_force[3576] <= 1'h0;
      write_done_data_log_force[3577] <= 1'h0;
      write_done_data_log_force[3578] <= 1'h0;
      write_done_data_log_force[3579] <= 1'h0;
      write_done_data_log_force[3580] <= 1'h0;
      write_done_data_log_force[3581] <= 1'h0;
      write_done_data_log_force[3582] <= 1'h0;
      write_done_data_log_force[3583] <= 1'h0;
      write_done_data_log_force[3584] <= 1'h0;
      write_done_data_log_force[3585] <= 1'h0;
      write_done_data_log_force[3586] <= 1'h0;
      write_done_data_log_force[3587] <= 1'h0;
      write_done_data_log_force[3588] <= 1'h0;
      write_done_data_log_force[3589] <= 1'h0;
      write_done_data_log_force[3590] <= 1'h0;
      write_done_data_log_force[3591] <= 1'h0;
      write_done_data_log_force[3592] <= 1'h0;
      write_done_data_log_force[3593] <= 1'h0;
      write_done_data_log_force[3594] <= 1'h0;
      write_done_data_log_force[3595] <= 1'h0;
      write_done_data_log_force[3596] <= 1'h0;
      write_done_data_log_force[3597] <= 1'h0;
      write_done_data_log_force[3598] <= 1'h0;
      write_done_data_log_force[3599] <= 1'h0;
      write_done_data_log_force[3600] <= 1'h0;
      write_done_data_log_force[3601] <= 1'h0;
      write_done_data_log_force[3602] <= 1'h0;
      write_done_data_log_force[3603] <= 1'h0;
      write_done_data_log_force[3604] <= 1'h0;
      write_done_data_log_force[3605] <= 1'h0;
      write_done_data_log_force[3606] <= 1'h0;
      write_done_data_log_force[3607] <= 1'h0;
      write_done_data_log_force[3608] <= 1'h0;
      write_done_data_log_force[3609] <= 1'h0;
      write_done_data_log_force[3610] <= 1'h0;
      write_done_data_log_force[3611] <= 1'h0;
      write_done_data_log_force[3612] <= 1'h0;
      write_done_data_log_force[3613] <= 1'h0;
      write_done_data_log_force[3614] <= 1'h0;
      write_done_data_log_force[3615] <= 1'h0;
      write_done_data_log_force[3616] <= 1'h0;
      write_done_data_log_force[3617] <= 1'h0;
      write_done_data_log_force[3618] <= 1'h0;
      write_done_data_log_force[3619] <= 1'h0;
      write_done_data_log_force[3620] <= 1'h0;
      write_done_data_log_force[3621] <= 1'h0;
      write_done_data_log_force[3622] <= 1'h0;
      write_done_data_log_force[3623] <= 1'h0;
      write_done_data_log_force[3624] <= 1'h0;
      write_done_data_log_force[3625] <= 1'h0;
      write_done_data_log_force[3626] <= 1'h0;
      write_done_data_log_force[3627] <= 1'h0;
      write_done_data_log_force[3628] <= 1'h0;
      write_done_data_log_force[3629] <= 1'h0;
      write_done_data_log_force[3630] <= 1'h0;
      write_done_data_log_force[3631] <= 1'h0;
      write_done_data_log_force[3632] <= 1'h0;
      write_done_data_log_force[3633] <= 1'h0;
      write_done_data_log_force[3634] <= 1'h0;
      write_done_data_log_force[3635] <= 1'h0;
      write_done_data_log_force[3636] <= 1'h0;
      write_done_data_log_force[3637] <= 1'h0;
      write_done_data_log_force[3638] <= 1'h0;
      write_done_data_log_force[3639] <= 1'h0;
      write_done_data_log_force[3640] <= 1'h0;
      write_done_data_log_force[3641] <= 1'h0;
      write_done_data_log_force[3642] <= 1'h0;
      write_done_data_log_force[3643] <= 1'h0;
      write_done_data_log_force[3644] <= 1'h0;
      write_done_data_log_force[3645] <= 1'h0;
      write_done_data_log_force[3646] <= 1'h0;
      write_done_data_log_force[3647] <= 1'h0;
      write_done_data_log_force[3648] <= 1'h0;
      write_done_data_log_force[3649] <= 1'h0;
      write_done_data_log_force[3650] <= 1'h0;
      write_done_data_log_force[3651] <= 1'h0;
      write_done_data_log_force[3652] <= 1'h0;
      write_done_data_log_force[3653] <= 1'h0;
      write_done_data_log_force[3654] <= 1'h0;
      write_done_data_log_force[3655] <= 1'h0;
      write_done_data_log_force[3656] <= 1'h0;
      write_done_data_log_force[3657] <= 1'h0;
      write_done_data_log_force[3658] <= 1'h0;
      write_done_data_log_force[3659] <= 1'h0;
      write_done_data_log_force[3660] <= 1'h0;
      write_done_data_log_force[3661] <= 1'h0;
      write_done_data_log_force[3662] <= 1'h0;
      write_done_data_log_force[3663] <= 1'h0;
      write_done_data_log_force[3664] <= 1'h0;
      write_done_data_log_force[3665] <= 1'h0;
      write_done_data_log_force[3666] <= 1'h0;
      write_done_data_log_force[3667] <= 1'h0;
      write_done_data_log_force[3668] <= 1'h0;
      write_done_data_log_force[3669] <= 1'h0;
      write_done_data_log_force[3670] <= 1'h0;
      write_done_data_log_force[3671] <= 1'h0;
      write_done_data_log_force[3672] <= 1'h0;
      write_done_data_log_force[3673] <= 1'h0;
      write_done_data_log_force[3674] <= 1'h0;
      write_done_data_log_force[3675] <= 1'h0;
      write_done_data_log_force[3676] <= 1'h0;
      write_done_data_log_force[3677] <= 1'h0;
      write_done_data_log_force[3678] <= 1'h0;
      write_done_data_log_force[3679] <= 1'h0;
      write_done_data_log_force[3680] <= 1'h0;
      write_done_data_log_force[3681] <= 1'h0;
      write_done_data_log_force[3682] <= 1'h0;
      write_done_data_log_force[3683] <= 1'h0;
      write_done_data_log_force[3684] <= 1'h0;
      write_done_data_log_force[3685] <= 1'h0;
      write_done_data_log_force[3686] <= 1'h0;
      write_done_data_log_force[3687] <= 1'h0;
      write_done_data_log_force[3688] <= 1'h0;
      write_done_data_log_force[3689] <= 1'h0;
      write_done_data_log_force[3690] <= 1'h0;
      write_done_data_log_force[3691] <= 1'h0;
      write_done_data_log_force[3692] <= 1'h0;
      write_done_data_log_force[3693] <= 1'h0;
      write_done_data_log_force[3694] <= 1'h0;
      write_done_data_log_force[3695] <= 1'h0;
      write_done_data_log_force[3696] <= 1'h0;
      write_done_data_log_force[3697] <= 1'h0;
      write_done_data_log_force[3698] <= 1'h0;
      write_done_data_log_force[3699] <= 1'h0;
      write_done_data_log_force[3700] <= 1'h0;
      write_done_data_log_force[3701] <= 1'h0;
      write_done_data_log_force[3702] <= 1'h0;
      write_done_data_log_force[3703] <= 1'h0;
      write_done_data_log_force[3704] <= 1'h0;
      write_done_data_log_force[3705] <= 1'h0;
      write_done_data_log_force[3706] <= 1'h0;
      write_done_data_log_force[3707] <= 1'h0;
      write_done_data_log_force[3708] <= 1'h0;
      write_done_data_log_force[3709] <= 1'h0;
      write_done_data_log_force[3710] <= 1'h0;
      write_done_data_log_force[3711] <= 1'h0;
      write_done_data_log_force[3712] <= 1'h0;
      write_done_data_log_force[3713] <= 1'h0;
      write_done_data_log_force[3714] <= 1'h0;
      write_done_data_log_force[3715] <= 1'h0;
      write_done_data_log_force[3716] <= 1'h0;
      write_done_data_log_force[3717] <= 1'h0;
      write_done_data_log_force[3718] <= 1'h0;
      write_done_data_log_force[3719] <= 1'h0;
      write_done_data_log_force[3720] <= 1'h0;
      write_done_data_log_force[3721] <= 1'h0;
      write_done_data_log_force[3722] <= 1'h0;
      write_done_data_log_force[3723] <= 1'h0;
      write_done_data_log_force[3724] <= 1'h0;
      write_done_data_log_force[3725] <= 1'h0;
      write_done_data_log_force[3726] <= 1'h0;
      write_done_data_log_force[3727] <= 1'h0;
      write_done_data_log_force[3728] <= 1'h0;
      write_done_data_log_force[3729] <= 1'h0;
      write_done_data_log_force[3730] <= 1'h0;
      write_done_data_log_force[3731] <= 1'h0;
      write_done_data_log_force[3732] <= 1'h0;
      write_done_data_log_force[3733] <= 1'h0;
      write_done_data_log_force[3734] <= 1'h0;
      write_done_data_log_force[3735] <= 1'h0;
      write_done_data_log_force[3736] <= 1'h0;
      write_done_data_log_force[3737] <= 1'h0;
      write_done_data_log_force[3738] <= 1'h0;
      write_done_data_log_force[3739] <= 1'h0;
      write_done_data_log_force[3740] <= 1'h0;
      write_done_data_log_force[3741] <= 1'h0;
      write_done_data_log_force[3742] <= 1'h0;
      write_done_data_log_force[3743] <= 1'h0;
      write_done_data_log_force[3744] <= 1'h0;
      write_done_data_log_force[3745] <= 1'h0;
      write_done_data_log_force[3746] <= 1'h0;
      write_done_data_log_force[3747] <= 1'h0;
      write_done_data_log_force[3748] <= 1'h0;
      write_done_data_log_force[3749] <= 1'h0;
      write_done_data_log_force[3750] <= 1'h0;
      write_done_data_log_force[3751] <= 1'h0;
      write_done_data_log_force[3752] <= 1'h0;
      write_done_data_log_force[3753] <= 1'h0;
      write_done_data_log_force[3754] <= 1'h0;
      write_done_data_log_force[3755] <= 1'h0;
      write_done_data_log_force[3756] <= 1'h0;
      write_done_data_log_force[3757] <= 1'h0;
      write_done_data_log_force[3758] <= 1'h0;
      write_done_data_log_force[3759] <= 1'h0;
      write_done_data_log_force[3760] <= 1'h0;
      write_done_data_log_force[3761] <= 1'h0;
      write_done_data_log_force[3762] <= 1'h0;
      write_done_data_log_force[3763] <= 1'h0;
      write_done_data_log_force[3764] <= 1'h0;
      write_done_data_log_force[3765] <= 1'h0;
      write_done_data_log_force[3766] <= 1'h0;
      write_done_data_log_force[3767] <= 1'h0;
      write_done_data_log_force[3768] <= 1'h0;
      write_done_data_log_force[3769] <= 1'h0;
      write_done_data_log_force[3770] <= 1'h0;
      write_done_data_log_force[3771] <= 1'h0;
      write_done_data_log_force[3772] <= 1'h0;
      write_done_data_log_force[3773] <= 1'h0;
      write_done_data_log_force[3774] <= 1'h0;
      write_done_data_log_force[3775] <= 1'h0;
      write_done_data_log_force[3776] <= 1'h0;
      write_done_data_log_force[3777] <= 1'h0;
      write_done_data_log_force[3778] <= 1'h0;
      write_done_data_log_force[3779] <= 1'h0;
      write_done_data_log_force[3780] <= 1'h0;
      write_done_data_log_force[3781] <= 1'h0;
      write_done_data_log_force[3782] <= 1'h0;
      write_done_data_log_force[3783] <= 1'h0;
      write_done_data_log_force[3784] <= 1'h0;
      write_done_data_log_force[3785] <= 1'h0;
      write_done_data_log_force[3786] <= 1'h0;
      write_done_data_log_force[3787] <= 1'h0;
      write_done_data_log_force[3788] <= 1'h0;
      write_done_data_log_force[3789] <= 1'h0;
      write_done_data_log_force[3790] <= 1'h0;
      write_done_data_log_force[3791] <= 1'h0;
      write_done_data_log_force[3792] <= 1'h0;
      write_done_data_log_force[3793] <= 1'h0;
      write_done_data_log_force[3794] <= 1'h0;
      write_done_data_log_force[3795] <= 1'h0;
      write_done_data_log_force[3796] <= 1'h0;
      write_done_data_log_force[3797] <= 1'h0;
      write_done_data_log_force[3798] <= 1'h0;
      write_done_data_log_force[3799] <= 1'h0;
      write_done_data_log_force[3800] <= 1'h0;
      write_done_data_log_force[3801] <= 1'h0;
      write_done_data_log_force[3802] <= 1'h0;
      write_done_data_log_force[3803] <= 1'h0;
      write_done_data_log_force[3804] <= 1'h0;
      write_done_data_log_force[3805] <= 1'h0;
      write_done_data_log_force[3806] <= 1'h0;
      write_done_data_log_force[3807] <= 1'h0;
      write_done_data_log_force[3808] <= 1'h0;
      write_done_data_log_force[3809] <= 1'h0;
      write_done_data_log_force[3810] <= 1'h0;
      write_done_data_log_force[3811] <= 1'h0;
      write_done_data_log_force[3812] <= 1'h0;
      write_done_data_log_force[3813] <= 1'h0;
      write_done_data_log_force[3814] <= 1'h0;
      write_done_data_log_force[3815] <= 1'h0;
      write_done_data_log_force[3816] <= 1'h0;
      write_done_data_log_force[3817] <= 1'h0;
      write_done_data_log_force[3818] <= 1'h0;
      write_done_data_log_force[3819] <= 1'h0;
      write_done_data_log_force[3820] <= 1'h0;
      write_done_data_log_force[3821] <= 1'h0;
      write_done_data_log_force[3822] <= 1'h0;
      write_done_data_log_force[3823] <= 1'h0;
      write_done_data_log_force[3824] <= 1'h0;
      write_done_data_log_force[3825] <= 1'h0;
      write_done_data_log_force[3826] <= 1'h0;
      write_done_data_log_force[3827] <= 1'h0;
      write_done_data_log_force[3828] <= 1'h0;
      write_done_data_log_force[3829] <= 1'h0;
      write_done_data_log_force[3830] <= 1'h0;
      write_done_data_log_force[3831] <= 1'h0;
      write_done_data_log_force[3832] <= 1'h0;
      write_done_data_log_force[3833] <= 1'h0;
      write_done_data_log_force[3834] <= 1'h0;
      write_done_data_log_force[3835] <= 1'h0;
      write_done_data_log_force[3836] <= 1'h0;
      write_done_data_log_force[3837] <= 1'h0;
      write_done_data_log_force[3838] <= 1'h0;
      write_done_data_log_force[3839] <= 1'h0;
      write_done_data_log_force[3840] <= 1'h0;
      write_done_data_log_force[3841] <= 1'h0;
      write_done_data_log_force[3842] <= 1'h0;
      write_done_data_log_force[3843] <= 1'h0;
      write_done_data_log_force[3844] <= 1'h0;
      write_done_data_log_force[3845] <= 1'h0;
      write_done_data_log_force[3846] <= 1'h0;
      write_done_data_log_force[3847] <= 1'h0;
      write_done_data_log_force[3848] <= 1'h0;
      write_done_data_log_force[3849] <= 1'h0;
      write_done_data_log_force[3850] <= 1'h0;
      write_done_data_log_force[3851] <= 1'h0;
      write_done_data_log_force[3852] <= 1'h0;
      write_done_data_log_force[3853] <= 1'h0;
      write_done_data_log_force[3854] <= 1'h0;
      write_done_data_log_force[3855] <= 1'h0;
      write_done_data_log_force[3856] <= 1'h0;
      write_done_data_log_force[3857] <= 1'h0;
      write_done_data_log_force[3858] <= 1'h0;
      write_done_data_log_force[3859] <= 1'h0;
      write_done_data_log_force[3860] <= 1'h0;
      write_done_data_log_force[3861] <= 1'h0;
      write_done_data_log_force[3862] <= 1'h0;
      write_done_data_log_force[3863] <= 1'h0;
      write_done_data_log_force[3864] <= 1'h0;
      write_done_data_log_force[3865] <= 1'h0;
      write_done_data_log_force[3866] <= 1'h0;
      write_done_data_log_force[3867] <= 1'h0;
      write_done_data_log_force[3868] <= 1'h0;
      write_done_data_log_force[3869] <= 1'h0;
      write_done_data_log_force[3870] <= 1'h0;
      write_done_data_log_force[3871] <= 1'h0;
      write_done_data_log_force[3872] <= 1'h0;
      write_done_data_log_force[3873] <= 1'h0;
      write_done_data_log_force[3874] <= 1'h0;
      write_done_data_log_force[3875] <= 1'h0;
      write_done_data_log_force[3876] <= 1'h0;
      write_done_data_log_force[3877] <= 1'h0;
      write_done_data_log_force[3878] <= 1'h0;
      write_done_data_log_force[3879] <= 1'h0;
      write_done_data_log_force[3880] <= 1'h0;
      write_done_data_log_force[3881] <= 1'h0;
      write_done_data_log_force[3882] <= 1'h0;
      write_done_data_log_force[3883] <= 1'h0;
      write_done_data_log_force[3884] <= 1'h0;
      write_done_data_log_force[3885] <= 1'h0;
      write_done_data_log_force[3886] <= 1'h0;
      write_done_data_log_force[3887] <= 1'h0;
      write_done_data_log_force[3888] <= 1'h0;
      write_done_data_log_force[3889] <= 1'h0;
      write_done_data_log_force[3890] <= 1'h0;
      write_done_data_log_force[3891] <= 1'h0;
      write_done_data_log_force[3892] <= 1'h0;
      write_done_data_log_force[3893] <= 1'h0;
      write_done_data_log_force[3894] <= 1'h0;
      write_done_data_log_force[3895] <= 1'h0;
      write_done_data_log_force[3896] <= 1'h0;
      write_done_data_log_force[3897] <= 1'h0;
      write_done_data_log_force[3898] <= 1'h0;
      write_done_data_log_force[3899] <= 1'h0;
      write_done_data_log_force[3900] <= 1'h0;
      write_done_data_log_force[3901] <= 1'h0;
      write_done_data_log_force[3902] <= 1'h0;
      write_done_data_log_force[3903] <= 1'h0;
      write_done_data_log_force[3904] <= 1'h0;
      write_done_data_log_force[3905] <= 1'h0;
      write_done_data_log_force[3906] <= 1'h0;
      write_done_data_log_force[3907] <= 1'h0;
      write_done_data_log_force[3908] <= 1'h0;
      write_done_data_log_force[3909] <= 1'h0;
      write_done_data_log_force[3910] <= 1'h0;
      write_done_data_log_force[3911] <= 1'h0;
      write_done_data_log_force[3912] <= 1'h0;
      write_done_data_log_force[3913] <= 1'h0;
      write_done_data_log_force[3914] <= 1'h0;
      write_done_data_log_force[3915] <= 1'h0;
      write_done_data_log_force[3916] <= 1'h0;
      write_done_data_log_force[3917] <= 1'h0;
      write_done_data_log_force[3918] <= 1'h0;
      write_done_data_log_force[3919] <= 1'h0;
      write_done_data_log_force[3920] <= 1'h0;
      write_done_data_log_force[3921] <= 1'h0;
      write_done_data_log_force[3922] <= 1'h0;
      write_done_data_log_force[3923] <= 1'h0;
      write_done_data_log_force[3924] <= 1'h0;
      write_done_data_log_force[3925] <= 1'h0;
      write_done_data_log_force[3926] <= 1'h0;
      write_done_data_log_force[3927] <= 1'h0;
      write_done_data_log_force[3928] <= 1'h0;
      write_done_data_log_force[3929] <= 1'h0;
      write_done_data_log_force[3930] <= 1'h0;
      write_done_data_log_force[3931] <= 1'h0;
      write_done_data_log_force[3932] <= 1'h0;
      write_done_data_log_force[3933] <= 1'h0;
      write_done_data_log_force[3934] <= 1'h0;
      write_done_data_log_force[3935] <= 1'h0;
      write_done_data_log_force[3936] <= 1'h0;
      write_done_data_log_force[3937] <= 1'h0;
      write_done_data_log_force[3938] <= 1'h0;
      write_done_data_log_force[3939] <= 1'h0;
      write_done_data_log_force[3940] <= 1'h0;
      write_done_data_log_force[3941] <= 1'h0;
      write_done_data_log_force[3942] <= 1'h0;
      write_done_data_log_force[3943] <= 1'h0;
      write_done_data_log_force[3944] <= 1'h0;
      write_done_data_log_force[3945] <= 1'h0;
      write_done_data_log_force[3946] <= 1'h0;
      write_done_data_log_force[3947] <= 1'h0;
      write_done_data_log_force[3948] <= 1'h0;
      write_done_data_log_force[3949] <= 1'h0;
      write_done_data_log_force[3950] <= 1'h0;
      write_done_data_log_force[3951] <= 1'h0;
      write_done_data_log_force[3952] <= 1'h0;
      write_done_data_log_force[3953] <= 1'h0;
      write_done_data_log_force[3954] <= 1'h0;
      write_done_data_log_force[3955] <= 1'h0;
      write_done_data_log_force[3956] <= 1'h0;
      write_done_data_log_force[3957] <= 1'h0;
      write_done_data_log_force[3958] <= 1'h0;
      write_done_data_log_force[3959] <= 1'h0;
      write_done_data_log_force[3960] <= 1'h0;
      write_done_data_log_force[3961] <= 1'h0;
      write_done_data_log_force[3962] <= 1'h0;
      write_done_data_log_force[3963] <= 1'h0;
      write_done_data_log_force[3964] <= 1'h0;
      write_done_data_log_force[3965] <= 1'h0;
      write_done_data_log_force[3966] <= 1'h0;
      write_done_data_log_force[3967] <= 1'h0;
      write_done_data_log_force[3968] <= 1'h0;
      write_done_data_log_force[3969] <= 1'h0;
      write_done_data_log_force[3970] <= 1'h0;
      write_done_data_log_force[3971] <= 1'h0;
      write_done_data_log_force[3972] <= 1'h0;
      write_done_data_log_force[3973] <= 1'h0;
      write_done_data_log_force[3974] <= 1'h0;
      write_done_data_log_force[3975] <= 1'h0;
      write_done_data_log_force[3976] <= 1'h0;
      write_done_data_log_force[3977] <= 1'h0;
      write_done_data_log_force[3978] <= 1'h0;
      write_done_data_log_force[3979] <= 1'h0;
      write_done_data_log_force[3980] <= 1'h0;
      write_done_data_log_force[3981] <= 1'h0;
      write_done_data_log_force[3982] <= 1'h0;
      write_done_data_log_force[3983] <= 1'h0;
      write_done_data_log_force[3984] <= 1'h0;
      write_done_data_log_force[3985] <= 1'h0;
      write_done_data_log_force[3986] <= 1'h0;
      write_done_data_log_force[3987] <= 1'h0;
      write_done_data_log_force[3988] <= 1'h0;
      write_done_data_log_force[3989] <= 1'h0;
      write_done_data_log_force[3990] <= 1'h0;
      write_done_data_log_force[3991] <= 1'h0;
      write_done_data_log_force[3992] <= 1'h0;
      write_done_data_log_force[3993] <= 1'h0;
      write_done_data_log_force[3994] <= 1'h0;
      write_done_data_log_force[3995] <= 1'h0;
      write_done_data_log_force[3996] <= 1'h0;
      write_done_data_log_force[3997] <= 1'h0;
      write_done_data_log_force[3998] <= 1'h0;
      write_done_data_log_force[3999] <= 1'h0;
      write_done_data_log_force[4000] <= 1'h0;
      write_done_data_log_force[4001] <= 1'h0;
      write_done_data_log_force[4002] <= 1'h0;
      write_done_data_log_force[4003] <= 1'h0;
      write_done_data_log_force[4004] <= 1'h0;
      write_done_data_log_force[4005] <= 1'h0;
      write_done_data_log_force[4006] <= 1'h0;
      write_done_data_log_force[4007] <= 1'h0;
      write_done_data_log_force[4008] <= 1'h0;
      write_done_data_log_force[4009] <= 1'h0;
      write_done_data_log_force[4010] <= 1'h0;
      write_done_data_log_force[4011] <= 1'h0;
      write_done_data_log_force[4012] <= 1'h0;
      write_done_data_log_force[4013] <= 1'h0;
      write_done_data_log_force[4014] <= 1'h0;
      write_done_data_log_force[4015] <= 1'h0;
      write_done_data_log_force[4016] <= 1'h0;
      write_done_data_log_force[4017] <= 1'h0;
      write_done_data_log_force[4018] <= 1'h0;
      write_done_data_log_force[4019] <= 1'h0;
      write_done_data_log_force[4020] <= 1'h0;
      write_done_data_log_force[4021] <= 1'h0;
      write_done_data_log_force[4022] <= 1'h0;
      write_done_data_log_force[4023] <= 1'h0;
      write_done_data_log_force[4024] <= 1'h0;
      write_done_data_log_force[4025] <= 1'h0;
      write_done_data_log_force[4026] <= 1'h0;
      write_done_data_log_force[4027] <= 1'h0;
      write_done_data_log_force[4028] <= 1'h0;
      write_done_data_log_force[4029] <= 1'h0;
      write_done_data_log_force[4030] <= 1'h0;
      write_done_data_log_force[4031] <= 1'h0;
      write_done_data_log_force[4032] <= 1'h0;
      write_done_data_log_force[4033] <= 1'h0;
      write_done_data_log_force[4034] <= 1'h0;
      write_done_data_log_force[4035] <= 1'h0;
      write_done_data_log_force[4036] <= 1'h0;
      write_done_data_log_force[4037] <= 1'h0;
      write_done_data_log_force[4038] <= 1'h0;
      write_done_data_log_force[4039] <= 1'h0;
      write_done_data_log_force[4040] <= 1'h0;
      write_done_data_log_force[4041] <= 1'h0;
      write_done_data_log_force[4042] <= 1'h0;
      write_done_data_log_force[4043] <= 1'h0;
      write_done_data_log_force[4044] <= 1'h0;
      write_done_data_log_force[4045] <= 1'h0;
      write_done_data_log_force[4046] <= 1'h0;
      write_done_data_log_force[4047] <= 1'h0;
      write_done_data_log_force[4048] <= 1'h0;
      write_done_data_log_force[4049] <= 1'h0;
      write_done_data_log_force[4050] <= 1'h0;
      write_done_data_log_force[4051] <= 1'h0;
      write_done_data_log_force[4052] <= 1'h0;
      write_done_data_log_force[4053] <= 1'h0;
      write_done_data_log_force[4054] <= 1'h0;
      write_done_data_log_force[4055] <= 1'h0;
      write_done_data_log_force[4056] <= 1'h0;
      write_done_data_log_force[4057] <= 1'h0;
      write_done_data_log_force[4058] <= 1'h0;
      write_done_data_log_force[4059] <= 1'h0;
      write_done_data_log_force[4060] <= 1'h0;
      write_done_data_log_force[4061] <= 1'h0;
      write_done_data_log_force[4062] <= 1'h0;
      write_done_data_log_force[4063] <= 1'h0;
      write_done_data_log_force[4064] <= 1'h0;
      write_done_data_log_force[4065] <= 1'h0;
      write_done_data_log_force[4066] <= 1'h0;
      write_done_data_log_force[4067] <= 1'h0;
      write_done_data_log_force[4068] <= 1'h0;
      write_done_data_log_force[4069] <= 1'h0;
      write_done_data_log_force[4070] <= 1'h0;
      write_done_data_log_force[4071] <= 1'h0;
      write_done_data_log_force[4072] <= 1'h0;
      write_done_data_log_force[4073] <= 1'h0;
      write_done_data_log_force[4074] <= 1'h0;
      write_done_data_log_force[4075] <= 1'h0;
      write_done_data_log_force[4076] <= 1'h0;
      write_done_data_log_force[4077] <= 1'h0;
      write_done_data_log_force[4078] <= 1'h0;
      write_done_data_log_force[4079] <= 1'h0;
      write_done_data_log_force[4080] <= 1'h0;
      write_done_data_log_force[4081] <= 1'h0;
      write_done_data_log_force[4082] <= 1'h0;
      write_done_data_log_force[4083] <= 1'h0;
      write_done_data_log_force[4084] <= 1'h0;
      write_done_data_log_force[4085] <= 1'h0;
      write_done_data_log_force[4086] <= 1'h0;
      write_done_data_log_force[4087] <= 1'h0;
      write_done_data_log_force[4088] <= 1'h0;
      write_done_data_log_force[4089] <= 1'h0;
      write_done_data_log_force[4090] <= 1'h0;
      write_done_data_log_force[4091] <= 1'h0;
      write_done_data_log_force[4092] <= 1'h0;
      write_done_data_log_force[4093] <= 1'h0;
      write_done_data_log_force[4094] <= 1'h0;
      write_done_data_log_force[4095] <= 1'h0;
      write_done_data_log_force[4096] <= 1'h0;
      write_done_data_log_force[4097] <= 1'h0;
      write_done_data_log_force[4098] <= 1'h0;
      write_done_data_log_force[4099] <= 1'h0;
      write_done_data_log_force[4100] <= 1'h0;
      write_done_data_log_force[4101] <= 1'h0;
      write_done_data_log_force[4102] <= 1'h0;
      write_done_data_log_force[4103] <= 1'h0;
      write_done_data_log_force[4104] <= 1'h0;
      write_done_data_log_force[4105] <= 1'h0;
      write_done_data_log_force[4106] <= 1'h0;
      write_done_data_log_force[4107] <= 1'h0;
      write_done_data_log_force[4108] <= 1'h0;
      write_done_data_log_force[4109] <= 1'h0;
      write_done_data_log_force[4110] <= 1'h0;
      write_done_data_log_force[4111] <= 1'h0;
      write_done_data_log_force[4112] <= 1'h0;
      write_done_data_log_force[4113] <= 1'h0;
      write_done_data_log_force[4114] <= 1'h0;
      write_done_data_log_force[4115] <= 1'h0;
      write_done_data_log_force[4116] <= 1'h0;
      write_done_data_log_force[4117] <= 1'h0;
      write_done_data_log_force[4118] <= 1'h0;
      write_done_data_log_force[4119] <= 1'h0;
      write_done_data_log_force[4120] <= 1'h0;
      write_done_data_log_force[4121] <= 1'h0;
      write_done_data_log_force[4122] <= 1'h0;
      write_done_data_log_force[4123] <= 1'h0;
      write_done_data_log_force[4124] <= 1'h0;
      write_done_data_log_force[4125] <= 1'h0;
      write_done_data_log_force[4126] <= 1'h0;
      write_done_data_log_force[4127] <= 1'h0;
      write_done_data_log_force[4128] <= 1'h0;
      write_done_data_log_force[4129] <= 1'h0;
      write_done_data_log_force[4130] <= 1'h0;
      write_done_data_log_force[4131] <= 1'h0;
      write_done_data_log_force[4132] <= 1'h0;
      write_done_data_log_force[4133] <= 1'h0;
      write_done_data_log_force[4134] <= 1'h0;
      write_done_data_log_force[4135] <= 1'h0;
      write_done_data_log_force[4136] <= 1'h0;
      write_done_data_log_force[4137] <= 1'h0;
      write_done_data_log_force[4138] <= 1'h0;
      write_done_data_log_force[4139] <= 1'h0;
      write_done_data_log_force[4140] <= 1'h0;
      write_done_data_log_force[4141] <= 1'h0;
      write_done_data_log_force[4142] <= 1'h0;
      write_done_data_log_force[4143] <= 1'h0;
      write_done_data_log_force[4144] <= 1'h0;
      write_done_data_log_force[4145] <= 1'h0;
      write_done_data_log_force[4146] <= 1'h0;
      write_done_data_log_force[4147] <= 1'h0;
      write_done_data_log_force[4148] <= 1'h0;
      write_done_data_log_force[4149] <= 1'h0;
      write_done_data_log_force[4150] <= 1'h0;
      write_done_data_log_force[4151] <= 1'h0;
      write_done_data_log_force[4152] <= 1'h0;
      write_done_data_log_force[4153] <= 1'h0;
      write_done_data_log_force[4154] <= 1'h0;
      write_done_data_log_force[4155] <= 1'h0;
      write_done_data_log_force[4156] <= 1'h0;
      write_done_data_log_force[4157] <= 1'h0;
      write_done_data_log_force[4158] <= 1'h0;
      write_done_data_log_force[4159] <= 1'h0;
      write_done_data_log_force[4160] <= 1'h0;
      write_done_data_log_force[4161] <= 1'h0;
      write_done_data_log_force[4162] <= 1'h0;
      write_done_data_log_force[4163] <= 1'h0;
      write_done_data_log_force[4164] <= 1'h0;
      write_done_data_log_force[4165] <= 1'h0;
      write_done_data_log_force[4166] <= 1'h0;
      write_done_data_log_force[4167] <= 1'h0;
      write_done_data_log_force[4168] <= 1'h0;
      write_done_data_log_force[4169] <= 1'h0;
      write_done_data_log_force[4170] <= 1'h0;
      write_done_data_log_force[4171] <= 1'h0;
      write_done_data_log_force[4172] <= 1'h0;
      write_done_data_log_force[4173] <= 1'h0;
      write_done_data_log_force[4174] <= 1'h0;
      write_done_data_log_force[4175] <= 1'h0;
      write_done_data_log_force[4176] <= 1'h0;
      write_done_data_log_force[4177] <= 1'h0;
      write_done_data_log_force[4178] <= 1'h0;
      write_done_data_log_force[4179] <= 1'h0;
      write_done_data_log_force[4180] <= 1'h0;
      write_done_data_log_force[4181] <= 1'h0;
      write_done_data_log_force[4182] <= 1'h0;
      write_done_data_log_force[4183] <= 1'h0;
      write_done_data_log_force[4184] <= 1'h0;
      write_done_data_log_force[4185] <= 1'h0;
      write_done_data_log_force[4186] <= 1'h0;
      write_done_data_log_force[4187] <= 1'h0;
      write_done_data_log_force[4188] <= 1'h0;
      write_done_data_log_force[4189] <= 1'h0;
      write_done_data_log_force[4190] <= 1'h0;
      write_done_data_log_force[4191] <= 1'h0;
      write_done_data_log_force[4192] <= 1'h0;
      write_done_data_log_force[4193] <= 1'h0;
      write_done_data_log_force[4194] <= 1'h0;
      write_done_data_log_force[4195] <= 1'h0;
      write_done_data_log_force[4196] <= 1'h0;
      write_done_data_log_force[4197] <= 1'h0;
      write_done_data_log_force[4198] <= 1'h0;
      write_done_data_log_force[4199] <= 1'h0;
      write_done_data_log_force[4200] <= 1'h0;
      write_done_data_log_force[4201] <= 1'h0;
      write_done_data_log_force[4202] <= 1'h0;
      write_done_data_log_force[4203] <= 1'h0;
      write_done_data_log_force[4204] <= 1'h0;
      write_done_data_log_force[4205] <= 1'h0;
      write_done_data_log_force[4206] <= 1'h0;
      write_done_data_log_force[4207] <= 1'h0;
      write_done_data_log_force[4208] <= 1'h0;
      write_done_data_log_force[4209] <= 1'h0;
      write_done_data_log_force[4210] <= 1'h0;
      write_done_data_log_force[4211] <= 1'h0;
      write_done_data_log_force[4212] <= 1'h0;
      write_done_data_log_force[4213] <= 1'h0;
      write_done_data_log_force[4214] <= 1'h0;
      write_done_data_log_force[4215] <= 1'h0;
      write_done_data_log_force[4216] <= 1'h0;
      write_done_data_log_force[4217] <= 1'h0;
      write_done_data_log_force[4218] <= 1'h0;
      write_done_data_log_force[4219] <= 1'h0;
      write_done_data_log_force[4220] <= 1'h0;
      write_done_data_log_force[4221] <= 1'h0;
      write_done_data_log_force[4222] <= 1'h0;
      write_done_data_log_force[4223] <= 1'h0;
      write_done_data_log_force[4224] <= 1'h0;
      write_done_data_log_force[4225] <= 1'h0;
      write_done_data_log_force[4226] <= 1'h0;
      write_done_data_log_force[4227] <= 1'h0;
      write_done_data_log_force[4228] <= 1'h0;
      write_done_data_log_force[4229] <= 1'h0;
      write_done_data_log_force[4230] <= 1'h0;
      write_done_data_log_force[4231] <= 1'h0;
      write_done_data_log_force[4232] <= 1'h0;
      write_done_data_log_force[4233] <= 1'h0;
      write_done_data_log_force[4234] <= 1'h0;
      write_done_data_log_force[4235] <= 1'h0;
      write_done_data_log_force[4236] <= 1'h0;
      write_done_data_log_force[4237] <= 1'h0;
      write_done_data_log_force[4238] <= 1'h0;
      write_done_data_log_force[4239] <= 1'h0;
      write_done_data_log_force[4240] <= 1'h0;
      write_done_data_log_force[4241] <= 1'h0;
      write_done_data_log_force[4242] <= 1'h0;
      write_done_data_log_force[4243] <= 1'h0;
      write_done_data_log_force[4244] <= 1'h0;
      write_done_data_log_force[4245] <= 1'h0;
      write_done_data_log_force[4246] <= 1'h0;
      write_done_data_log_force[4247] <= 1'h0;
      write_done_data_log_force[4248] <= 1'h0;
      write_done_data_log_force[4249] <= 1'h0;
      write_done_data_log_force[4250] <= 1'h0;
      write_done_data_log_force[4251] <= 1'h0;
      write_done_data_log_force[4252] <= 1'h0;
      write_done_data_log_force[4253] <= 1'h0;
      write_done_data_log_force[4254] <= 1'h0;
      write_done_data_log_force[4255] <= 1'h0;
      write_done_data_log_force[4256] <= 1'h0;
      write_done_data_log_force[4257] <= 1'h0;
      write_done_data_log_force[4258] <= 1'h0;
      write_done_data_log_force[4259] <= 1'h0;
      write_done_data_log_force[4260] <= 1'h0;
      write_done_data_log_force[4261] <= 1'h0;
      write_done_data_log_force[4262] <= 1'h0;
      write_done_data_log_force[4263] <= 1'h0;
      write_done_data_log_force[4264] <= 1'h0;
      write_done_data_log_force[4265] <= 1'h0;
      write_done_data_log_force[4266] <= 1'h0;
      write_done_data_log_force[4267] <= 1'h0;
      write_done_data_log_force[4268] <= 1'h0;
      write_done_data_log_force[4269] <= 1'h0;
      write_done_data_log_force[4270] <= 1'h0;
      write_done_data_log_force[4271] <= 1'h0;
      write_done_data_log_force[4272] <= 1'h0;
      write_done_data_log_force[4273] <= 1'h0;
      write_done_data_log_force[4274] <= 1'h0;
      write_done_data_log_force[4275] <= 1'h0;
      write_done_data_log_force[4276] <= 1'h0;
      write_done_data_log_force[4277] <= 1'h0;
      write_done_data_log_force[4278] <= 1'h0;
      write_done_data_log_force[4279] <= 1'h0;
      write_done_data_log_force[4280] <= 1'h0;
      write_done_data_log_force[4281] <= 1'h0;
      write_done_data_log_force[4282] <= 1'h0;
      write_done_data_log_force[4283] <= 1'h0;
      write_done_data_log_force[4284] <= 1'h0;
      write_done_data_log_force[4285] <= 1'h0;
      write_done_data_log_force[4286] <= 1'h0;
      write_done_data_log_force[4287] <= 1'h0;
      write_done_data_log_force[4288] <= 1'h0;
      write_done_data_log_force[4289] <= 1'h0;
      write_done_data_log_force[4290] <= 1'h0;
      write_done_data_log_force[4291] <= 1'h0;
      write_done_data_log_force[4292] <= 1'h0;
      write_done_data_log_force[4293] <= 1'h0;
      write_done_data_log_force[4294] <= 1'h0;
      write_done_data_log_force[4295] <= 1'h0;
      write_done_data_log_force[4296] <= 1'h0;
      write_done_data_log_force[4297] <= 1'h0;
      write_done_data_log_force[4298] <= 1'h0;
      write_done_data_log_force[4299] <= 1'h0;
      write_done_data_log_force[4300] <= 1'h0;
      write_done_data_log_force[4301] <= 1'h0;
      write_done_data_log_force[4302] <= 1'h0;
      write_done_data_log_force[4303] <= 1'h0;
      write_done_data_log_force[4304] <= 1'h0;
      write_done_data_log_force[4305] <= 1'h0;
      write_done_data_log_force[4306] <= 1'h0;
      write_done_data_log_force[4307] <= 1'h0;
      write_done_data_log_force[4308] <= 1'h0;
      write_done_data_log_force[4309] <= 1'h0;
      write_done_data_log_force[4310] <= 1'h0;
      write_done_data_log_force[4311] <= 1'h0;
      write_done_data_log_force[4312] <= 1'h0;
      write_done_data_log_force[4313] <= 1'h0;
      write_done_data_log_force[4314] <= 1'h0;
      write_done_data_log_force[4315] <= 1'h0;
      write_done_data_log_force[4316] <= 1'h0;
      write_done_data_log_force[4317] <= 1'h0;
      write_done_data_log_force[4318] <= 1'h0;
      write_done_data_log_force[4319] <= 1'h0;
      write_done_data_log_force[4320] <= 1'h0;
      write_done_data_log_force[4321] <= 1'h0;
      write_done_data_log_force[4322] <= 1'h0;
      write_done_data_log_force[4323] <= 1'h0;
      write_done_data_log_force[4324] <= 1'h0;
      write_done_data_log_force[4325] <= 1'h0;
      write_done_data_log_force[4326] <= 1'h0;
      write_done_data_log_force[4327] <= 1'h0;
      write_done_data_log_force[4328] <= 1'h0;
      write_done_data_log_force[4329] <= 1'h0;
      write_done_data_log_force[4330] <= 1'h0;
      write_done_data_log_force[4331] <= 1'h0;
      write_done_data_log_force[4332] <= 1'h0;
      write_done_data_log_force[4333] <= 1'h0;
      write_done_data_log_force[4334] <= 1'h0;
      write_done_data_log_force[4335] <= 1'h0;
      write_done_data_log_force[4336] <= 1'h0;
      write_done_data_log_force[4337] <= 1'h0;
      write_done_data_log_force[4338] <= 1'h0;
      write_done_data_log_force[4339] <= 1'h0;
      write_done_data_log_force[4340] <= 1'h0;
      write_done_data_log_force[4341] <= 1'h0;
      write_done_data_log_force[4342] <= 1'h0;
      write_done_data_log_force[4343] <= 1'h0;
      write_done_data_log_force[4344] <= 1'h0;
      write_done_data_log_force[4345] <= 1'h0;
      write_done_data_log_force[4346] <= 1'h0;
      write_done_data_log_force[4347] <= 1'h0;
      write_done_data_log_force[4348] <= 1'h0;
      write_done_data_log_force[4349] <= 1'h0;
      write_done_data_log_force[4350] <= 1'h0;
      write_done_data_log_force[4351] <= 1'h0;
      write_done_data_log_force[4352] <= 1'h0;
      write_done_data_log_force[4353] <= 1'h0;
      write_done_data_log_force[4354] <= 1'h0;
      write_done_data_log_force[4355] <= 1'h0;
      write_done_data_log_force[4356] <= 1'h0;
      write_done_data_log_force[4357] <= 1'h0;
      write_done_data_log_force[4358] <= 1'h0;
      write_done_data_log_force[4359] <= 1'h0;
      write_done_data_log_force[4360] <= 1'h0;
      write_done_data_log_force[4361] <= 1'h0;
      write_done_data_log_force[4362] <= 1'h0;
      write_done_data_log_force[4363] <= 1'h0;
      write_done_data_log_force[4364] <= 1'h0;
      write_done_data_log_force[4365] <= 1'h0;
      write_done_data_log_force[4366] <= 1'h0;
      write_done_data_log_force[4367] <= 1'h0;
      write_done_data_log_force[4368] <= 1'h0;
      write_done_data_log_force[4369] <= 1'h0;
      write_done_data_log_force[4370] <= 1'h0;
      write_done_data_log_force[4371] <= 1'h0;
      write_done_data_log_force[4372] <= 1'h0;
      write_done_data_log_force[4373] <= 1'h0;
      write_done_data_log_force[4374] <= 1'h0;
      write_done_data_log_force[4375] <= 1'h0;
      write_done_data_log_force[4376] <= 1'h0;
      write_done_data_log_force[4377] <= 1'h0;
      write_done_data_log_force[4378] <= 1'h0;
      write_done_data_log_force[4379] <= 1'h0;
      write_done_data_log_force[4380] <= 1'h0;
      write_done_data_log_force[4381] <= 1'h0;
      write_done_data_log_force[4382] <= 1'h0;
      write_done_data_log_force[4383] <= 1'h0;
      write_done_data_log_force[4384] <= 1'h0;
      write_done_data_log_force[4385] <= 1'h0;
      write_done_data_log_force[4386] <= 1'h0;
      write_done_data_log_force[4387] <= 1'h0;
      write_done_data_log_force[4388] <= 1'h0;
      write_done_data_log_force[4389] <= 1'h0;
      write_done_data_log_force[4390] <= 1'h0;
      write_done_data_log_force[4391] <= 1'h0;
      write_done_data_log_force[4392] <= 1'h0;
      write_done_data_log_force[4393] <= 1'h0;
      write_done_data_log_force[4394] <= 1'h0;
      write_done_data_log_force[4395] <= 1'h0;
      write_done_data_log_force[4396] <= 1'h0;
      write_done_data_log_force[4397] <= 1'h0;
      write_done_data_log_force[4398] <= 1'h0;
      write_done_data_log_force[4399] <= 1'h0;
      write_done_data_log_force[4400] <= 1'h0;
      write_done_data_log_force[4401] <= 1'h0;
      write_done_data_log_force[4402] <= 1'h0;
      write_done_data_log_force[4403] <= 1'h0;
      write_done_data_log_force[4404] <= 1'h0;
      write_done_data_log_force[4405] <= 1'h0;
      write_done_data_log_force[4406] <= 1'h0;
      write_done_data_log_force[4407] <= 1'h0;
      write_done_data_log_force[4408] <= 1'h0;
      write_done_data_log_force[4409] <= 1'h0;
      write_done_data_log_force[4410] <= 1'h0;
      write_done_data_log_force[4411] <= 1'h0;
      write_done_data_log_force[4412] <= 1'h0;
      write_done_data_log_force[4413] <= 1'h0;
      write_done_data_log_force[4414] <= 1'h0;
      write_done_data_log_force[4415] <= 1'h0;
      write_done_data_log_force[4416] <= 1'h0;
      write_done_data_log_force[4417] <= 1'h0;
      write_done_data_log_force[4418] <= 1'h0;
      write_done_data_log_force[4419] <= 1'h0;
      write_done_data_log_force[4420] <= 1'h0;
      write_done_data_log_force[4421] <= 1'h0;
      write_done_data_log_force[4422] <= 1'h0;
      write_done_data_log_force[4423] <= 1'h0;
      write_done_data_log_force[4424] <= 1'h0;
      write_done_data_log_force[4425] <= 1'h0;
      write_done_data_log_force[4426] <= 1'h0;
      write_done_data_log_force[4427] <= 1'h0;
      write_done_data_log_force[4428] <= 1'h0;
      write_done_data_log_force[4429] <= 1'h0;
      write_done_data_log_force[4430] <= 1'h0;
      write_done_data_log_force[4431] <= 1'h0;
      write_done_data_log_force[4432] <= 1'h0;
      write_done_data_log_force[4433] <= 1'h0;
      write_done_data_log_force[4434] <= 1'h0;
      write_done_data_log_force[4435] <= 1'h0;
      write_done_data_log_force[4436] <= 1'h0;
      write_done_data_log_force[4437] <= 1'h0;
      write_done_data_log_force[4438] <= 1'h0;
      write_done_data_log_force[4439] <= 1'h0;
      write_done_data_log_force[4440] <= 1'h0;
      write_done_data_log_force[4441] <= 1'h0;
      write_done_data_log_force[4442] <= 1'h0;
      write_done_data_log_force[4443] <= 1'h0;
      write_done_data_log_force[4444] <= 1'h0;
      write_done_data_log_force[4445] <= 1'h0;
      write_done_data_log_force[4446] <= 1'h0;
      write_done_data_log_force[4447] <= 1'h0;
      write_done_data_log_force[4448] <= 1'h0;
      write_done_data_log_force[4449] <= 1'h0;
      write_done_data_log_force[4450] <= 1'h0;
      write_done_data_log_force[4451] <= 1'h0;
      write_done_data_log_force[4452] <= 1'h0;
      write_done_data_log_force[4453] <= 1'h0;
      write_done_data_log_force[4454] <= 1'h0;
      write_done_data_log_force[4455] <= 1'h0;
      write_done_data_log_force[4456] <= 1'h0;
      write_done_data_log_force[4457] <= 1'h0;
      write_done_data_log_force[4458] <= 1'h0;
      write_done_data_log_force[4459] <= 1'h0;
      write_done_data_log_force[4460] <= 1'h0;
      write_done_data_log_force[4461] <= 1'h0;
      write_done_data_log_force[4462] <= 1'h0;
      write_done_data_log_force[4463] <= 1'h0;
      write_done_data_log_force[4464] <= 1'h0;
      write_done_data_log_force[4465] <= 1'h0;
      write_done_data_log_force[4466] <= 1'h0;
      write_done_data_log_force[4467] <= 1'h0;
      write_done_data_log_force[4468] <= 1'h0;
      write_done_data_log_force[4469] <= 1'h0;
      write_done_data_log_force[4470] <= 1'h0;
      write_done_data_log_force[4471] <= 1'h0;
      write_done_data_log_force[4472] <= 1'h0;
      write_done_data_log_force[4473] <= 1'h0;
      write_done_data_log_force[4474] <= 1'h0;
      write_done_data_log_force[4475] <= 1'h0;
      write_done_data_log_force[4476] <= 1'h0;
      write_done_data_log_force[4477] <= 1'h0;
      write_done_data_log_force[4478] <= 1'h0;
      write_done_data_log_force[4479] <= 1'h0;
      write_done_data_log_force[4480] <= 1'h0;
      write_done_data_log_force[4481] <= 1'h0;
      write_done_data_log_force[4482] <= 1'h0;
      write_done_data_log_force[4483] <= 1'h0;
      write_done_data_log_force[4484] <= 1'h0;
      write_done_data_log_force[4485] <= 1'h0;
      write_done_data_log_force[4486] <= 1'h0;
      write_done_data_log_force[4487] <= 1'h0;
      write_done_data_log_force[4488] <= 1'h0;
      write_done_data_log_force[4489] <= 1'h0;
      write_done_data_log_force[4490] <= 1'h0;
      write_done_data_log_force[4491] <= 1'h0;
      write_done_data_log_force[4492] <= 1'h0;
      write_done_data_log_force[4493] <= 1'h0;
      write_done_data_log_force[4494] <= 1'h0;
      write_done_data_log_force[4495] <= 1'h0;
      write_done_data_log_force[4496] <= 1'h0;
      write_done_data_log_force[4497] <= 1'h0;
      write_done_data_log_force[4498] <= 1'h0;
      write_done_data_log_force[4499] <= 1'h0;
      write_done_data_log_force[4500] <= 1'h0;
      write_done_data_log_force[4501] <= 1'h0;
      write_done_data_log_force[4502] <= 1'h0;
      write_done_data_log_force[4503] <= 1'h0;
      write_done_data_log_force[4504] <= 1'h0;
      write_done_data_log_force[4505] <= 1'h0;
      write_done_data_log_force[4506] <= 1'h0;
      write_done_data_log_force[4507] <= 1'h0;
      write_done_data_log_force[4508] <= 1'h0;
      write_done_data_log_force[4509] <= 1'h0;
      write_done_data_log_force[4510] <= 1'h0;
      write_done_data_log_force[4511] <= 1'h0;
      write_done_data_log_force[4512] <= 1'h0;
      write_done_data_log_force[4513] <= 1'h0;
      write_done_data_log_force[4514] <= 1'h0;
      write_done_data_log_force[4515] <= 1'h0;
      write_done_data_log_force[4516] <= 1'h0;
      write_done_data_log_force[4517] <= 1'h0;
      write_done_data_log_force[4518] <= 1'h0;
      write_done_data_log_force[4519] <= 1'h0;
      write_done_data_log_force[4520] <= 1'h0;
      write_done_data_log_force[4521] <= 1'h0;
      write_done_data_log_force[4522] <= 1'h0;
      write_done_data_log_force[4523] <= 1'h0;
      write_done_data_log_force[4524] <= 1'h0;
      write_done_data_log_force[4525] <= 1'h0;
      write_done_data_log_force[4526] <= 1'h0;
      write_done_data_log_force[4527] <= 1'h0;
      write_done_data_log_force[4528] <= 1'h0;
      write_done_data_log_force[4529] <= 1'h0;
      write_done_data_log_force[4530] <= 1'h0;
      write_done_data_log_force[4531] <= 1'h0;
      write_done_data_log_force[4532] <= 1'h0;
      write_done_data_log_force[4533] <= 1'h0;
      write_done_data_log_force[4534] <= 1'h0;
      write_done_data_log_force[4535] <= 1'h0;
      write_done_data_log_force[4536] <= 1'h0;
      write_done_data_log_force[4537] <= 1'h0;
      write_done_data_log_force[4538] <= 1'h0;
      write_done_data_log_force[4539] <= 1'h0;
      write_done_data_log_force[4540] <= 1'h0;
      write_done_data_log_force[4541] <= 1'h0;
      write_done_data_log_force[4542] <= 1'h0;
      write_done_data_log_force[4543] <= 1'h0;
      write_done_data_log_force[4544] <= 1'h0;
      write_done_data_log_force[4545] <= 1'h0;
      write_done_data_log_force[4546] <= 1'h0;
      write_done_data_log_force[4547] <= 1'h0;
      write_done_data_log_force[4548] <= 1'h0;
      write_done_data_log_force[4549] <= 1'h0;
      write_done_data_log_force[4550] <= 1'h0;
      write_done_data_log_force[4551] <= 1'h0;
      write_done_data_log_force[4552] <= 1'h0;
      write_done_data_log_force[4553] <= 1'h0;
      write_done_data_log_force[4554] <= 1'h0;
      write_done_data_log_force[4555] <= 1'h0;
      write_done_data_log_force[4556] <= 1'h0;
      write_done_data_log_force[4557] <= 1'h0;
      write_done_data_log_force[4558] <= 1'h0;
      write_done_data_log_force[4559] <= 1'h0;
      write_done_data_log_force[4560] <= 1'h0;
      write_done_data_log_force[4561] <= 1'h0;
      write_done_data_log_force[4562] <= 1'h0;
      write_done_data_log_force[4563] <= 1'h0;
      write_done_data_log_force[4564] <= 1'h0;
      write_done_data_log_force[4565] <= 1'h0;
      write_done_data_log_force[4566] <= 1'h0;
      write_done_data_log_force[4567] <= 1'h0;
      write_done_data_log_force[4568] <= 1'h0;
      write_done_data_log_force[4569] <= 1'h0;
      write_done_data_log_force[4570] <= 1'h0;
      write_done_data_log_force[4571] <= 1'h0;
      write_done_data_log_force[4572] <= 1'h0;
      write_done_data_log_force[4573] <= 1'h0;
      write_done_data_log_force[4574] <= 1'h0;
      write_done_data_log_force[4575] <= 1'h0;
      write_done_data_log_force[4576] <= 1'h0;
      write_done_data_log_force[4577] <= 1'h0;
      write_done_data_log_force[4578] <= 1'h0;
      write_done_data_log_force[4579] <= 1'h0;
      write_done_data_log_force[4580] <= 1'h0;
      write_done_data_log_force[4581] <= 1'h0;
      write_done_data_log_force[4582] <= 1'h0;
      write_done_data_log_force[4583] <= 1'h0;
      write_done_data_log_force[4584] <= 1'h0;
      write_done_data_log_force[4585] <= 1'h0;
      write_done_data_log_force[4586] <= 1'h0;
      write_done_data_log_force[4587] <= 1'h0;
      write_done_data_log_force[4588] <= 1'h0;
      write_done_data_log_force[4589] <= 1'h0;
      write_done_data_log_force[4590] <= 1'h0;
      write_done_data_log_force[4591] <= 1'h0;
      write_done_data_log_force[4592] <= 1'h0;
      write_done_data_log_force[4593] <= 1'h0;
      write_done_data_log_force[4594] <= 1'h0;
      write_done_data_log_force[4595] <= 1'h0;
      write_done_data_log_force[4596] <= 1'h0;
      write_done_data_log_force[4597] <= 1'h0;
      write_done_data_log_force[4598] <= 1'h0;
      write_done_data_log_force[4599] <= 1'h0;
      write_done_data_log_force[4600] <= 1'h0;
      write_done_data_log_force[4601] <= 1'h0;
      write_done_data_log_force[4602] <= 1'h0;
      write_done_data_log_force[4603] <= 1'h0;
      write_done_data_log_force[4604] <= 1'h0;
      write_done_data_log_force[4605] <= 1'h0;
      write_done_data_log_force[4606] <= 1'h0;
      write_done_data_log_force[4607] <= 1'h0;
      write_done_data_log_force[4608] <= 1'h0;
      write_done_data_log_force[4609] <= 1'h0;
      write_done_data_log_force[4610] <= 1'h0;
      write_done_data_log_force[4611] <= 1'h0;
      write_done_data_log_force[4612] <= 1'h0;
      write_done_data_log_force[4613] <= 1'h0;
      write_done_data_log_force[4614] <= 1'h0;
      write_done_data_log_force[4615] <= 1'h0;
      write_done_data_log_force[4616] <= 1'h0;
      write_done_data_log_force[4617] <= 1'h0;
      write_done_data_log_force[4618] <= 1'h0;
      write_done_data_log_force[4619] <= 1'h0;
      write_done_data_log_force[4620] <= 1'h0;
      write_done_data_log_force[4621] <= 1'h0;
      write_done_data_log_force[4622] <= 1'h0;
      write_done_data_log_force[4623] <= 1'h0;
      write_done_data_log_force[4624] <= 1'h0;
      write_done_data_log_force[4625] <= 1'h0;
      write_done_data_log_force[4626] <= 1'h0;
      write_done_data_log_force[4627] <= 1'h0;
      write_done_data_log_force[4628] <= 1'h0;
      write_done_data_log_force[4629] <= 1'h0;
      write_done_data_log_force[4630] <= 1'h0;
      write_done_data_log_force[4631] <= 1'h0;
      write_done_data_log_force[4632] <= 1'h0;
      write_done_data_log_force[4633] <= 1'h0;
      write_done_data_log_force[4634] <= 1'h0;
      write_done_data_log_force[4635] <= 1'h0;
      write_done_data_log_force[4636] <= 1'h0;
      write_done_data_log_force[4637] <= 1'h0;
      write_done_data_log_force[4638] <= 1'h0;
      write_done_data_log_force[4639] <= 1'h0;
      write_done_data_log_force[4640] <= 1'h0;
      write_done_data_log_force[4641] <= 1'h0;
      write_done_data_log_force[4642] <= 1'h0;
      write_done_data_log_force[4643] <= 1'h0;
      write_done_data_log_force[4644] <= 1'h0;
      write_done_data_log_force[4645] <= 1'h0;
      write_done_data_log_force[4646] <= 1'h0;
      write_done_data_log_force[4647] <= 1'h0;
      write_done_data_log_force[4648] <= 1'h0;
      write_done_data_log_force[4649] <= 1'h0;
      write_done_data_log_force[4650] <= 1'h0;
      write_done_data_log_force[4651] <= 1'h0;
      write_done_data_log_force[4652] <= 1'h0;
      write_done_data_log_force[4653] <= 1'h0;
      write_done_data_log_force[4654] <= 1'h0;
      write_done_data_log_force[4655] <= 1'h0;
      write_done_data_log_force[4656] <= 1'h0;
      write_done_data_log_force[4657] <= 1'h0;
      write_done_data_log_force[4658] <= 1'h0;
      write_done_data_log_force[4659] <= 1'h0;
      write_done_data_log_force[4660] <= 1'h0;
      write_done_data_log_force[4661] <= 1'h0;
      write_done_data_log_force[4662] <= 1'h0;
      write_done_data_log_force[4663] <= 1'h0;
      write_done_data_log_force[4664] <= 1'h0;
      write_done_data_log_force[4665] <= 1'h0;
      write_done_data_log_force[4666] <= 1'h0;
      write_done_data_log_force[4667] <= 1'h0;
      write_done_data_log_force[4668] <= 1'h0;
      write_done_data_log_force[4669] <= 1'h0;
      write_done_data_log_force[4670] <= 1'h0;
      write_done_data_log_force[4671] <= 1'h0;
      write_done_data_log_force[4672] <= 1'h0;
      write_done_data_log_force[4673] <= 1'h0;
      write_done_data_log_force[4674] <= 1'h0;
      write_done_data_log_force[4675] <= 1'h0;
      write_done_data_log_force[4676] <= 1'h0;
      write_done_data_log_force[4677] <= 1'h0;
      write_done_data_log_force[4678] <= 1'h0;
      write_done_data_log_force[4679] <= 1'h0;
      write_done_data_log_force[4680] <= 1'h0;
      write_done_data_log_force[4681] <= 1'h0;
      write_done_data_log_force[4682] <= 1'h0;
      write_done_data_log_force[4683] <= 1'h0;
      write_done_data_log_force[4684] <= 1'h0;
      write_done_data_log_force[4685] <= 1'h0;
      write_done_data_log_force[4686] <= 1'h0;
      write_done_data_log_force[4687] <= 1'h0;
      write_done_data_log_force[4688] <= 1'h0;
      write_done_data_log_force[4689] <= 1'h0;
      write_done_data_log_force[4690] <= 1'h0;
      write_done_data_log_force[4691] <= 1'h0;
      write_done_data_log_force[4692] <= 1'h0;
      write_done_data_log_force[4693] <= 1'h0;
      write_done_data_log_force[4694] <= 1'h0;
      write_done_data_log_force[4695] <= 1'h0;
      write_done_data_log_force[4696] <= 1'h0;
      write_done_data_log_force[4697] <= 1'h0;
      write_done_data_log_force[4698] <= 1'h0;
      write_done_data_log_force[4699] <= 1'h0;
      write_done_data_log_force[4700] <= 1'h0;
      write_done_data_log_force[4701] <= 1'h0;
      write_done_data_log_force[4702] <= 1'h0;
      write_done_data_log_force[4703] <= 1'h0;
      write_done_data_log_force[4704] <= 1'h0;
      write_done_data_log_force[4705] <= 1'h0;
      write_done_data_log_force[4706] <= 1'h0;
      write_done_data_log_force[4707] <= 1'h0;
      write_done_data_log_force[4708] <= 1'h0;
      write_done_data_log_force[4709] <= 1'h0;
      write_done_data_log_force[4710] <= 1'h0;
      write_done_data_log_force[4711] <= 1'h0;
      write_done_data_log_force[4712] <= 1'h0;
      write_done_data_log_force[4713] <= 1'h0;
      write_done_data_log_force[4714] <= 1'h0;
      write_done_data_log_force[4715] <= 1'h0;
      write_done_data_log_force[4716] <= 1'h0;
      write_done_data_log_force[4717] <= 1'h0;
      write_done_data_log_force[4718] <= 1'h0;
      write_done_data_log_force[4719] <= 1'h0;
      write_done_data_log_force[4720] <= 1'h0;
      write_done_data_log_force[4721] <= 1'h0;
      write_done_data_log_force[4722] <= 1'h0;
      write_done_data_log_force[4723] <= 1'h0;
      write_done_data_log_force[4724] <= 1'h0;
      write_done_data_log_force[4725] <= 1'h0;
      write_done_data_log_force[4726] <= 1'h0;
      write_done_data_log_force[4727] <= 1'h0;
      write_done_data_log_force[4728] <= 1'h0;
      write_done_data_log_force[4729] <= 1'h0;
      write_done_data_log_force[4730] <= 1'h0;
      write_done_data_log_force[4731] <= 1'h0;
      write_done_data_log_force[4732] <= 1'h0;
      write_done_data_log_force[4733] <= 1'h0;
      write_done_data_log_force[4734] <= 1'h0;
      write_done_data_log_force[4735] <= 1'h0;
      write_done_data_log_force[4736] <= 1'h0;
      write_done_data_log_force[4737] <= 1'h0;
      write_done_data_log_force[4738] <= 1'h0;
      write_done_data_log_force[4739] <= 1'h0;
      write_done_data_log_force[4740] <= 1'h0;
      write_done_data_log_force[4741] <= 1'h0;
      write_done_data_log_force[4742] <= 1'h0;
      write_done_data_log_force[4743] <= 1'h0;
      write_done_data_log_force[4744] <= 1'h0;
      write_done_data_log_force[4745] <= 1'h0;
      write_done_data_log_force[4746] <= 1'h0;
      write_done_data_log_force[4747] <= 1'h0;
      write_done_data_log_force[4748] <= 1'h0;
      write_done_data_log_force[4749] <= 1'h0;
      write_done_data_log_force[4750] <= 1'h0;
      write_done_data_log_force[4751] <= 1'h0;
      write_done_data_log_force[4752] <= 1'h0;
      write_done_data_log_force[4753] <= 1'h0;
      write_done_data_log_force[4754] <= 1'h0;
      write_done_data_log_force[4755] <= 1'h0;
      write_done_data_log_force[4756] <= 1'h0;
      write_done_data_log_force[4757] <= 1'h0;
      write_done_data_log_force[4758] <= 1'h0;
      write_done_data_log_force[4759] <= 1'h0;
      write_done_data_log_force[4760] <= 1'h0;
      write_done_data_log_force[4761] <= 1'h0;
      write_done_data_log_force[4762] <= 1'h0;
      write_done_data_log_force[4763] <= 1'h0;
      write_done_data_log_force[4764] <= 1'h0;
      write_done_data_log_force[4765] <= 1'h0;
      write_done_data_log_force[4766] <= 1'h0;
      write_done_data_log_force[4767] <= 1'h0;
      write_done_data_log_force[4768] <= 1'h0;
      write_done_data_log_force[4769] <= 1'h0;
      write_done_data_log_force[4770] <= 1'h0;
      write_done_data_log_force[4771] <= 1'h0;
      write_done_data_log_force[4772] <= 1'h0;
      write_done_data_log_force[4773] <= 1'h0;
      write_done_data_log_force[4774] <= 1'h0;
      write_done_data_log_force[4775] <= 1'h0;
      write_done_data_log_force[4776] <= 1'h0;
      write_done_data_log_force[4777] <= 1'h0;
      write_done_data_log_force[4778] <= 1'h0;
      write_done_data_log_force[4779] <= 1'h0;
      write_done_data_log_force[4780] <= 1'h0;
      write_done_data_log_force[4781] <= 1'h0;
      write_done_data_log_force[4782] <= 1'h0;
      write_done_data_log_force[4783] <= 1'h0;
      write_done_data_log_force[4784] <= 1'h0;
      write_done_data_log_force[4785] <= 1'h0;
      write_done_data_log_force[4786] <= 1'h0;
      write_done_data_log_force[4787] <= 1'h0;
      write_done_data_log_force[4788] <= 1'h0;
      write_done_data_log_force[4789] <= 1'h0;
      write_done_data_log_force[4790] <= 1'h0;
      write_done_data_log_force[4791] <= 1'h0;
      write_done_data_log_force[4792] <= 1'h0;
      write_done_data_log_force[4793] <= 1'h0;
      write_done_data_log_force[4794] <= 1'h0;
      write_done_data_log_force[4795] <= 1'h0;
      write_done_data_log_force[4796] <= 1'h0;
      write_done_data_log_force[4797] <= 1'h0;
      write_done_data_log_force[4798] <= 1'h0;
      write_done_data_log_force[4799] <= 1'h0;
      write_done_data_log_force[4800] <= 1'h0;
      write_done_data_log_force[4801] <= 1'h0;
      write_done_data_log_force[4802] <= 1'h0;
      write_done_data_log_force[4803] <= 1'h0;
      write_done_data_log_force[4804] <= 1'h0;
      write_done_data_log_force[4805] <= 1'h0;
      write_done_data_log_force[4806] <= 1'h0;
      write_done_data_log_force[4807] <= 1'h0;
      write_done_data_log_force[4808] <= 1'h0;
      write_done_data_log_force[4809] <= 1'h0;
      write_done_data_log_force[4810] <= 1'h0;
      write_done_data_log_force[4811] <= 1'h0;
      write_done_data_log_force[4812] <= 1'h0;
      write_done_data_log_force[4813] <= 1'h0;
      write_done_data_log_force[4814] <= 1'h0;
      write_done_data_log_force[4815] <= 1'h0;
      write_done_data_log_force[4816] <= 1'h0;
      write_done_data_log_force[4817] <= 1'h0;
      write_done_data_log_force[4818] <= 1'h0;
      write_done_data_log_force[4819] <= 1'h0;
      write_done_data_log_force[4820] <= 1'h0;
      write_done_data_log_force[4821] <= 1'h0;
      write_done_data_log_force[4822] <= 1'h0;
      write_done_data_log_force[4823] <= 1'h0;
      write_done_data_log_force[4824] <= 1'h0;
      write_done_data_log_force[4825] <= 1'h0;
      write_done_data_log_force[4826] <= 1'h0;
      write_done_data_log_force[4827] <= 1'h0;
      write_done_data_log_force[4828] <= 1'h0;
      write_done_data_log_force[4829] <= 1'h0;
      write_done_data_log_force[4830] <= 1'h0;
      write_done_data_log_force[4831] <= 1'h0;
      write_done_data_log_force[4832] <= 1'h0;
      write_done_data_log_force[4833] <= 1'h0;
      write_done_data_log_force[4834] <= 1'h0;
      write_done_data_log_force[4835] <= 1'h0;
      write_done_data_log_force[4836] <= 1'h0;
      write_done_data_log_force[4837] <= 1'h0;
      write_done_data_log_force[4838] <= 1'h0;
      write_done_data_log_force[4839] <= 1'h0;
      write_done_data_log_force[4840] <= 1'h0;
      write_done_data_log_force[4841] <= 1'h0;
      write_done_data_log_force[4842] <= 1'h0;
      write_done_data_log_force[4843] <= 1'h0;
      write_done_data_log_force[4844] <= 1'h0;
      write_done_data_log_force[4845] <= 1'h0;
      write_done_data_log_force[4846] <= 1'h0;
      write_done_data_log_force[4847] <= 1'h0;
      write_done_data_log_force[4848] <= 1'h0;
      write_done_data_log_force[4849] <= 1'h0;
      write_done_data_log_force[4850] <= 1'h0;
      write_done_data_log_force[4851] <= 1'h0;
      write_done_data_log_force[4852] <= 1'h0;
      write_done_data_log_force[4853] <= 1'h0;
      write_done_data_log_force[4854] <= 1'h0;
      write_done_data_log_force[4855] <= 1'h0;
      write_done_data_log_force[4856] <= 1'h0;
      write_done_data_log_force[4857] <= 1'h0;
      write_done_data_log_force[4858] <= 1'h0;
      write_done_data_log_force[4859] <= 1'h0;
      write_done_data_log_force[4860] <= 1'h0;
      write_done_data_log_force[4861] <= 1'h0;
      write_done_data_log_force[4862] <= 1'h0;
      write_done_data_log_force[4863] <= 1'h0;
      write_done_data_log_force[4864] <= 1'h0;
      write_done_data_log_force[4865] <= 1'h0;
      write_done_data_log_force[4866] <= 1'h0;
      write_done_data_log_force[4867] <= 1'h0;
      write_done_data_log_force[4868] <= 1'h0;
      write_done_data_log_force[4869] <= 1'h0;
      write_done_data_log_force[4870] <= 1'h0;
      write_done_data_log_force[4871] <= 1'h0;
      write_done_data_log_force[4872] <= 1'h0;
      write_done_data_log_force[4873] <= 1'h0;
      write_done_data_log_force[4874] <= 1'h0;
      write_done_data_log_force[4875] <= 1'h0;
      write_done_data_log_force[4876] <= 1'h0;
      write_done_data_log_force[4877] <= 1'h0;
      write_done_data_log_force[4878] <= 1'h0;
      write_done_data_log_force[4879] <= 1'h0;
      write_done_data_log_force[4880] <= 1'h0;
      write_done_data_log_force[4881] <= 1'h0;
      write_done_data_log_force[4882] <= 1'h0;
      write_done_data_log_force[4883] <= 1'h0;
      write_done_data_log_force[4884] <= 1'h0;
      write_done_data_log_force[4885] <= 1'h0;
      write_done_data_log_force[4886] <= 1'h0;
      write_done_data_log_force[4887] <= 1'h0;
      write_done_data_log_force[4888] <= 1'h0;
      write_done_data_log_force[4889] <= 1'h0;
      write_done_data_log_force[4890] <= 1'h0;
      write_done_data_log_force[4891] <= 1'h0;
      write_done_data_log_force[4892] <= 1'h0;
      write_done_data_log_force[4893] <= 1'h0;
      write_done_data_log_force[4894] <= 1'h0;
      write_done_data_log_force[4895] <= 1'h0;
      write_done_data_log_force[4896] <= 1'h0;
      write_done_data_log_force[4897] <= 1'h0;
      write_done_data_log_force[4898] <= 1'h0;
      write_done_data_log_force[4899] <= 1'h0;
      write_done_data_log_force[4900] <= 1'h0;
      write_done_data_log_force[4901] <= 1'h0;
      write_done_data_log_force[4902] <= 1'h0;
      write_done_data_log_force[4903] <= 1'h0;
      write_done_data_log_force[4904] <= 1'h0;
      write_done_data_log_force[4905] <= 1'h0;
      write_done_data_log_force[4906] <= 1'h0;
      write_done_data_log_force[4907] <= 1'h0;
      write_done_data_log_force[4908] <= 1'h0;
      write_done_data_log_force[4909] <= 1'h0;
      write_done_data_log_force[4910] <= 1'h0;
      write_done_data_log_force[4911] <= 1'h0;
      write_done_data_log_force[4912] <= 1'h0;
      write_done_data_log_force[4913] <= 1'h0;
      write_done_data_log_force[4914] <= 1'h0;
      write_done_data_log_force[4915] <= 1'h0;
      write_done_data_log_force[4916] <= 1'h0;
      write_done_data_log_force[4917] <= 1'h0;
      write_done_data_log_force[4918] <= 1'h0;
      write_done_data_log_force[4919] <= 1'h0;
      write_done_data_log_force[4920] <= 1'h0;
      write_done_data_log_force[4921] <= 1'h0;
      write_done_data_log_force[4922] <= 1'h0;
      write_done_data_log_force[4923] <= 1'h0;
      write_done_data_log_force[4924] <= 1'h0;
      write_done_data_log_force[4925] <= 1'h0;
      write_done_data_log_force[4926] <= 1'h0;
      write_done_data_log_force[4927] <= 1'h0;
      write_done_data_log_force[4928] <= 1'h0;
      write_done_data_log_force[4929] <= 1'h0;
      write_done_data_log_force[4930] <= 1'h0;
      write_done_data_log_force[4931] <= 1'h0;
      write_done_data_log_force[4932] <= 1'h0;
      write_done_data_log_force[4933] <= 1'h0;
      write_done_data_log_force[4934] <= 1'h0;
      write_done_data_log_force[4935] <= 1'h0;
      write_done_data_log_force[4936] <= 1'h0;
      write_done_data_log_force[4937] <= 1'h0;
      write_done_data_log_force[4938] <= 1'h0;
      write_done_data_log_force[4939] <= 1'h0;
      write_done_data_log_force[4940] <= 1'h0;
      write_done_data_log_force[4941] <= 1'h0;
      write_done_data_log_force[4942] <= 1'h0;
      write_done_data_log_force[4943] <= 1'h0;
      write_done_data_log_force[4944] <= 1'h0;
      write_done_data_log_force[4945] <= 1'h0;
      write_done_data_log_force[4946] <= 1'h0;
      write_done_data_log_force[4947] <= 1'h0;
      write_done_data_log_force[4948] <= 1'h0;
      write_done_data_log_force[4949] <= 1'h0;
      write_done_data_log_force[4950] <= 1'h0;
      write_done_data_log_force[4951] <= 1'h0;
      write_done_data_log_force[4952] <= 1'h0;
      write_done_data_log_force[4953] <= 1'h0;
      write_done_data_log_force[4954] <= 1'h0;
      write_done_data_log_force[4955] <= 1'h0;
      write_done_data_log_force[4956] <= 1'h0;
      write_done_data_log_force[4957] <= 1'h0;
      write_done_data_log_force[4958] <= 1'h0;
      write_done_data_log_force[4959] <= 1'h0;
      write_done_data_log_force[4960] <= 1'h0;
      write_done_data_log_force[4961] <= 1'h0;
      write_done_data_log_force[4962] <= 1'h0;
      write_done_data_log_force[4963] <= 1'h0;
      write_done_data_log_force[4964] <= 1'h0;
      write_done_data_log_force[4965] <= 1'h0;
      write_done_data_log_force[4966] <= 1'h0;
      write_done_data_log_force[4967] <= 1'h0;
      write_done_data_log_force[4968] <= 1'h0;
      write_done_data_log_force[4969] <= 1'h0;
      write_done_data_log_force[4970] <= 1'h0;
      write_done_data_log_force[4971] <= 1'h0;
      write_done_data_log_force[4972] <= 1'h0;
      write_done_data_log_force[4973] <= 1'h0;
      write_done_data_log_force[4974] <= 1'h0;
      write_done_data_log_force[4975] <= 1'h0;
      write_done_data_log_force[4976] <= 1'h0;
      write_done_data_log_force[4977] <= 1'h0;
      write_done_data_log_force[4978] <= 1'h0;
      write_done_data_log_force[4979] <= 1'h0;
      write_done_data_log_force[4980] <= 1'h0;
      write_done_data_log_force[4981] <= 1'h0;
      write_done_data_log_force[4982] <= 1'h0;
      write_done_data_log_force[4983] <= 1'h0;
      write_done_data_log_force[4984] <= 1'h0;
      write_done_data_log_force[4985] <= 1'h0;
      write_done_data_log_force[4986] <= 1'h0;
      write_done_data_log_force[4987] <= 1'h0;
      write_done_data_log_force[4988] <= 1'h0;
      write_done_data_log_force[4989] <= 1'h0;
      write_done_data_log_force[4990] <= 1'h0;
      write_done_data_log_force[4991] <= 1'h0;
      write_done_data_log_force[4992] <= 1'h0;
      write_done_data_log_force[4993] <= 1'h0;
      write_done_data_log_force[4994] <= 1'h0;
      write_done_data_log_force[4995] <= 1'h0;
      write_done_data_log_force[4996] <= 1'h0;
      write_done_data_log_force[4997] <= 1'h0;
      write_done_data_log_force[4998] <= 1'h0;
      write_done_data_log_force[4999] <= 1'h0;
      write_done_data_log_force[5000] <= 1'h0;
      write_done_data_log_force[5001] <= 1'h0;
      write_done_data_log_force[5002] <= 1'h0;
      write_done_data_log_force[5003] <= 1'h0;
      write_done_data_log_force[5004] <= 1'h0;
      write_done_data_log_force[5005] <= 1'h0;
      write_done_data_log_force[5006] <= 1'h0;
      write_done_data_log_force[5007] <= 1'h0;
      write_done_data_log_force[5008] <= 1'h0;
      write_done_data_log_force[5009] <= 1'h0;
      write_done_data_log_force[5010] <= 1'h0;
      write_done_data_log_force[5011] <= 1'h0;
      write_done_data_log_force[5012] <= 1'h0;
      write_done_data_log_force[5013] <= 1'h0;
      write_done_data_log_force[5014] <= 1'h0;
      write_done_data_log_force[5015] <= 1'h0;
      write_done_data_log_force[5016] <= 1'h0;
      write_done_data_log_force[5017] <= 1'h0;
      write_done_data_log_force[5018] <= 1'h0;
      write_done_data_log_force[5019] <= 1'h0;
      write_done_data_log_force[5020] <= 1'h0;
      write_done_data_log_force[5021] <= 1'h0;
      write_done_data_log_force[5022] <= 1'h0;
      write_done_data_log_force[5023] <= 1'h0;
      write_done_data_log_force[5024] <= 1'h0;
      write_done_data_log_force[5025] <= 1'h0;
      write_done_data_log_force[5026] <= 1'h0;
      write_done_data_log_force[5027] <= 1'h0;
      write_done_data_log_force[5028] <= 1'h0;
      write_done_data_log_force[5029] <= 1'h0;
      write_done_data_log_force[5030] <= 1'h0;
      write_done_data_log_force[5031] <= 1'h0;
      write_done_data_log_force[5032] <= 1'h0;
      write_done_data_log_force[5033] <= 1'h0;
      write_done_data_log_force[5034] <= 1'h0;
      write_done_data_log_force[5035] <= 1'h0;
      write_done_data_log_force[5036] <= 1'h0;
      write_done_data_log_force[5037] <= 1'h0;
      write_done_data_log_force[5038] <= 1'h0;
      write_done_data_log_force[5039] <= 1'h0;
      write_done_data_log_force[5040] <= 1'h0;
      write_done_data_log_force[5041] <= 1'h0;
      write_done_data_log_force[5042] <= 1'h0;
      write_done_data_log_force[5043] <= 1'h0;
      write_done_data_log_force[5044] <= 1'h0;
      write_done_data_log_force[5045] <= 1'h0;
      write_done_data_log_force[5046] <= 1'h0;
      write_done_data_log_force[5047] <= 1'h0;
      write_done_data_log_force[5048] <= 1'h0;
      write_done_data_log_force[5049] <= 1'h0;
      write_done_data_log_force[5050] <= 1'h0;
      write_done_data_log_force[5051] <= 1'h0;
      write_done_data_log_force[5052] <= 1'h0;
      write_done_data_log_force[5053] <= 1'h0;
      write_done_data_log_force[5054] <= 1'h0;
      write_done_data_log_force[5055] <= 1'h0;
      write_done_data_log_force[5056] <= 1'h0;
      write_done_data_log_force[5057] <= 1'h0;
      write_done_data_log_force[5058] <= 1'h0;
      write_done_data_log_force[5059] <= 1'h0;
      write_done_data_log_force[5060] <= 1'h0;
      write_done_data_log_force[5061] <= 1'h0;
      write_done_data_log_force[5062] <= 1'h0;
      write_done_data_log_force[5063] <= 1'h0;
      write_done_data_log_force[5064] <= 1'h0;
      write_done_data_log_force[5065] <= 1'h0;
      write_done_data_log_force[5066] <= 1'h0;
      write_done_data_log_force[5067] <= 1'h0;
      write_done_data_log_force[5068] <= 1'h0;
      write_done_data_log_force[5069] <= 1'h0;
      write_done_data_log_force[5070] <= 1'h0;
      write_done_data_log_force[5071] <= 1'h0;
      write_done_data_log_force[5072] <= 1'h0;
      write_done_data_log_force[5073] <= 1'h0;
      write_done_data_log_force[5074] <= 1'h0;
      write_done_data_log_force[5075] <= 1'h0;
      write_done_data_log_force[5076] <= 1'h0;
      write_done_data_log_force[5077] <= 1'h0;
      write_done_data_log_force[5078] <= 1'h0;
      write_done_data_log_force[5079] <= 1'h0;
      write_done_data_log_force[5080] <= 1'h0;
      write_done_data_log_force[5081] <= 1'h0;
      write_done_data_log_force[5082] <= 1'h0;
      write_done_data_log_force[5083] <= 1'h0;
      write_done_data_log_force[5084] <= 1'h0;
      write_done_data_log_force[5085] <= 1'h0;
      write_done_data_log_force[5086] <= 1'h0;
      write_done_data_log_force[5087] <= 1'h0;
      write_done_data_log_force[5088] <= 1'h0;
      write_done_data_log_force[5089] <= 1'h0;
      write_done_data_log_force[5090] <= 1'h0;
      write_done_data_log_force[5091] <= 1'h0;
      write_done_data_log_force[5092] <= 1'h0;
      write_done_data_log_force[5093] <= 1'h0;
      write_done_data_log_force[5094] <= 1'h0;
      write_done_data_log_force[5095] <= 1'h0;
      write_done_data_log_force[5096] <= 1'h0;
      write_done_data_log_force[5097] <= 1'h0;
      write_done_data_log_force[5098] <= 1'h0;
      write_done_data_log_force[5099] <= 1'h0;
      write_done_data_log_force[5100] <= 1'h0;
      write_done_data_log_force[5101] <= 1'h0;
      write_done_data_log_force[5102] <= 1'h0;
      write_done_data_log_force[5103] <= 1'h0;
      write_done_data_log_force[5104] <= 1'h0;
      write_done_data_log_force[5105] <= 1'h0;
      write_done_data_log_force[5106] <= 1'h0;
      write_done_data_log_force[5107] <= 1'h0;
      write_done_data_log_force[5108] <= 1'h0;
      write_done_data_log_force[5109] <= 1'h0;
      write_done_data_log_force[5110] <= 1'h0;
      write_done_data_log_force[5111] <= 1'h0;
      write_done_data_log_force[5112] <= 1'h0;
      write_done_data_log_force[5113] <= 1'h0;
      write_done_data_log_force[5114] <= 1'h0;
      write_done_data_log_force[5115] <= 1'h0;
      write_done_data_log_force[5116] <= 1'h0;
      write_done_data_log_force[5117] <= 1'h0;
      write_done_data_log_force[5118] <= 1'h0;
      write_done_data_log_force[5119] <= 1'h0;
      write_done_data_log_force[5120] <= 1'h0;
      write_done_data_log_force[5121] <= 1'h0;
      write_done_data_log_force[5122] <= 1'h0;
      write_done_data_log_force[5123] <= 1'h0;
      write_done_data_log_force[5124] <= 1'h0;
      write_done_data_log_force[5125] <= 1'h0;
      write_done_data_log_force[5126] <= 1'h0;
      write_done_data_log_force[5127] <= 1'h0;
      write_done_data_log_force[5128] <= 1'h0;
      write_done_data_log_force[5129] <= 1'h0;
      write_done_data_log_force[5130] <= 1'h0;
      write_done_data_log_force[5131] <= 1'h0;
      write_done_data_log_force[5132] <= 1'h0;
      write_done_data_log_force[5133] <= 1'h0;
      write_done_data_log_force[5134] <= 1'h0;
      write_done_data_log_force[5135] <= 1'h0;
      write_done_data_log_force[5136] <= 1'h0;
      write_done_data_log_force[5137] <= 1'h0;
      write_done_data_log_force[5138] <= 1'h0;
      write_done_data_log_force[5139] <= 1'h0;
      write_done_data_log_force[5140] <= 1'h0;
      write_done_data_log_force[5141] <= 1'h0;
      write_done_data_log_force[5142] <= 1'h0;
      write_done_data_log_force[5143] <= 1'h0;
      write_done_data_log_force[5144] <= 1'h0;
      write_done_data_log_force[5145] <= 1'h0;
      write_done_data_log_force[5146] <= 1'h0;
      write_done_data_log_force[5147] <= 1'h0;
      write_done_data_log_force[5148] <= 1'h0;
      write_done_data_log_force[5149] <= 1'h0;
      write_done_data_log_force[5150] <= 1'h0;
      write_done_data_log_force[5151] <= 1'h0;
      write_done_data_log_force[5152] <= 1'h0;
      write_done_data_log_force[5153] <= 1'h0;
      write_done_data_log_force[5154] <= 1'h0;
      write_done_data_log_force[5155] <= 1'h0;
      write_done_data_log_force[5156] <= 1'h0;
      write_done_data_log_force[5157] <= 1'h0;
      write_done_data_log_force[5158] <= 1'h0;
      write_done_data_log_force[5159] <= 1'h0;
      write_done_data_log_force[5160] <= 1'h0;
      write_done_data_log_force[5161] <= 1'h0;
      write_done_data_log_force[5162] <= 1'h0;
      write_done_data_log_force[5163] <= 1'h0;
      write_done_data_log_force[5164] <= 1'h0;
      write_done_data_log_force[5165] <= 1'h0;
      write_done_data_log_force[5166] <= 1'h0;
      write_done_data_log_force[5167] <= 1'h0;
      write_done_data_log_force[5168] <= 1'h0;
      write_done_data_log_force[5169] <= 1'h0;
      write_done_data_log_force[5170] <= 1'h0;
      write_done_data_log_force[5171] <= 1'h0;
      write_done_data_log_force[5172] <= 1'h0;
      write_done_data_log_force[5173] <= 1'h0;
      write_done_data_log_force[5174] <= 1'h0;
      write_done_data_log_force[5175] <= 1'h0;
      write_done_data_log_force[5176] <= 1'h0;
      write_done_data_log_force[5177] <= 1'h0;
      write_done_data_log_force[5178] <= 1'h0;
      write_done_data_log_force[5179] <= 1'h0;
      write_done_data_log_force[5180] <= 1'h0;
      write_done_data_log_force[5181] <= 1'h0;
      write_done_data_log_force[5182] <= 1'h0;
      write_done_data_log_force[5183] <= 1'h0;
      write_done_data_log_force[5184] <= 1'h0;
      write_done_data_log_force[5185] <= 1'h0;
      write_done_data_log_force[5186] <= 1'h0;
      write_done_data_log_force[5187] <= 1'h0;
      write_done_data_log_force[5188] <= 1'h0;
      write_done_data_log_force[5189] <= 1'h0;
      write_done_data_log_force[5190] <= 1'h0;
      write_done_data_log_force[5191] <= 1'h0;
      write_done_data_log_force[5192] <= 1'h0;
      write_done_data_log_force[5193] <= 1'h0;
      write_done_data_log_force[5194] <= 1'h0;
      write_done_data_log_force[5195] <= 1'h0;
      write_done_data_log_force[5196] <= 1'h0;
      write_done_data_log_force[5197] <= 1'h0;
      write_done_data_log_force[5198] <= 1'h0;
      write_done_data_log_force[5199] <= 1'h0;
      write_done_data_log_force[5200] <= 1'h0;
      write_done_data_log_force[5201] <= 1'h0;
      write_done_data_log_force[5202] <= 1'h0;
      write_done_data_log_force[5203] <= 1'h0;
      write_done_data_log_force[5204] <= 1'h0;
      write_done_data_log_force[5205] <= 1'h0;
      write_done_data_log_force[5206] <= 1'h0;
      write_done_data_log_force[5207] <= 1'h0;
      write_done_data_log_force[5208] <= 1'h0;
      write_done_data_log_force[5209] <= 1'h0;
      write_done_data_log_force[5210] <= 1'h0;
      write_done_data_log_force[5211] <= 1'h0;
      write_done_data_log_force[5212] <= 1'h0;
      write_done_data_log_force[5213] <= 1'h0;
      write_done_data_log_force[5214] <= 1'h0;
      write_done_data_log_force[5215] <= 1'h0;
      write_done_data_log_force[5216] <= 1'h0;
      write_done_data_log_force[5217] <= 1'h0;
      write_done_data_log_force[5218] <= 1'h0;
      write_done_data_log_force[5219] <= 1'h0;
      write_done_data_log_force[5220] <= 1'h0;
      write_done_data_log_force[5221] <= 1'h0;
      write_done_data_log_force[5222] <= 1'h0;
      write_done_data_log_force[5223] <= 1'h0;
      write_done_data_log_force[5224] <= 1'h0;
      write_done_data_log_force[5225] <= 1'h0;
      write_done_data_log_force[5226] <= 1'h0;
      write_done_data_log_force[5227] <= 1'h0;
      write_done_data_log_force[5228] <= 1'h0;
      write_done_data_log_force[5229] <= 1'h0;
      write_done_data_log_force[5230] <= 1'h0;
      write_done_data_log_force[5231] <= 1'h0;
      write_done_data_log_force[5232] <= 1'h0;
      write_done_data_log_force[5233] <= 1'h0;
      write_done_data_log_force[5234] <= 1'h0;
      write_done_data_log_force[5235] <= 1'h0;
      write_done_data_log_force[5236] <= 1'h0;
      write_done_data_log_force[5237] <= 1'h0;
      write_done_data_log_force[5238] <= 1'h0;
      write_done_data_log_force[5239] <= 1'h0;
      write_done_data_log_force[5240] <= 1'h0;
      write_done_data_log_force[5241] <= 1'h0;
      write_done_data_log_force[5242] <= 1'h0;
      write_done_data_log_force[5243] <= 1'h0;
      write_done_data_log_force[5244] <= 1'h0;
      write_done_data_log_force[5245] <= 1'h0;
      write_done_data_log_force[5246] <= 1'h0;
      write_done_data_log_force[5247] <= 1'h0;
      write_done_data_log_force[5248] <= 1'h0;
      write_done_data_log_force[5249] <= 1'h0;
      write_done_data_log_force[5250] <= 1'h0;
      write_done_data_log_force[5251] <= 1'h0;
      write_done_data_log_force[5252] <= 1'h0;
      write_done_data_log_force[5253] <= 1'h0;
      write_done_data_log_force[5254] <= 1'h0;
      write_done_data_log_force[5255] <= 1'h0;
      write_done_data_log_force[5256] <= 1'h0;
      write_done_data_log_force[5257] <= 1'h0;
      write_done_data_log_force[5258] <= 1'h0;
      write_done_data_log_force[5259] <= 1'h0;
      write_done_data_log_force[5260] <= 1'h0;
      write_done_data_log_force[5261] <= 1'h0;
      write_done_data_log_force[5262] <= 1'h0;
      write_done_data_log_force[5263] <= 1'h0;
      write_done_data_log_force[5264] <= 1'h0;
      write_done_data_log_force[5265] <= 1'h0;
      write_done_data_log_force[5266] <= 1'h0;
      write_done_data_log_force[5267] <= 1'h0;
      write_done_data_log_force[5268] <= 1'h0;
      write_done_data_log_force[5269] <= 1'h0;
      write_done_data_log_force[5270] <= 1'h0;
      write_done_data_log_force[5271] <= 1'h0;
      write_done_data_log_force[5272] <= 1'h0;
      write_done_data_log_force[5273] <= 1'h0;
      write_done_data_log_force[5274] <= 1'h0;
      write_done_data_log_force[5275] <= 1'h0;
      write_done_data_log_force[5276] <= 1'h0;
      write_done_data_log_force[5277] <= 1'h0;
      write_done_data_log_force[5278] <= 1'h0;
      write_done_data_log_force[5279] <= 1'h0;
      write_done_data_log_force[5280] <= 1'h0;
      write_done_data_log_force[5281] <= 1'h0;
      write_done_data_log_force[5282] <= 1'h0;
      write_done_data_log_force[5283] <= 1'h0;
      write_done_data_log_force[5284] <= 1'h0;
      write_done_data_log_force[5285] <= 1'h0;
      write_done_data_log_force[5286] <= 1'h0;
      write_done_data_log_force[5287] <= 1'h0;
      write_done_data_log_force[5288] <= 1'h0;
      write_done_data_log_force[5289] <= 1'h0;
      write_done_data_log_force[5290] <= 1'h0;
      write_done_data_log_force[5291] <= 1'h0;
      write_done_data_log_force[5292] <= 1'h0;
      write_done_data_log_force[5293] <= 1'h0;
      write_done_data_log_force[5294] <= 1'h0;
      write_done_data_log_force[5295] <= 1'h0;
      write_done_data_log_force[5296] <= 1'h0;
      write_done_data_log_force[5297] <= 1'h0;
      write_done_data_log_force[5298] <= 1'h0;
      write_done_data_log_force[5299] <= 1'h0;
      write_done_data_log_force[5300] <= 1'h0;
      write_done_data_log_force[5301] <= 1'h0;
      write_done_data_log_force[5302] <= 1'h0;
      write_done_data_log_force[5303] <= 1'h0;
      write_done_data_log_force[5304] <= 1'h0;
      write_done_data_log_force[5305] <= 1'h0;
      write_done_data_log_force[5306] <= 1'h0;
      write_done_data_log_force[5307] <= 1'h0;
      write_done_data_log_force[5308] <= 1'h0;
      write_done_data_log_force[5309] <= 1'h0;
      write_done_data_log_force[5310] <= 1'h0;
      write_done_data_log_force[5311] <= 1'h0;
      write_done_data_log_force[5312] <= 1'h0;
      write_done_data_log_force[5313] <= 1'h0;
      write_done_data_log_force[5314] <= 1'h0;
      write_done_data_log_force[5315] <= 1'h0;
      write_done_data_log_force[5316] <= 1'h0;
      write_done_data_log_force[5317] <= 1'h0;
      write_done_data_log_force[5318] <= 1'h0;
      write_done_data_log_force[5319] <= 1'h0;
      write_done_data_log_force[5320] <= 1'h0;
      write_done_data_log_force[5321] <= 1'h0;
      write_done_data_log_force[5322] <= 1'h0;
      write_done_data_log_force[5323] <= 1'h0;
      write_done_data_log_force[5324] <= 1'h0;
      write_done_data_log_force[5325] <= 1'h0;
      write_done_data_log_force[5326] <= 1'h0;
      write_done_data_log_force[5327] <= 1'h0;
      write_done_data_log_force[5328] <= 1'h0;
      write_done_data_log_force[5329] <= 1'h0;
      write_done_data_log_force[5330] <= 1'h0;
      write_done_data_log_force[5331] <= 1'h0;
      write_done_data_log_force[5332] <= 1'h0;
      write_done_data_log_force[5333] <= 1'h0;
      write_done_data_log_force[5334] <= 1'h0;
      write_done_data_log_force[5335] <= 1'h0;
      write_done_data_log_force[5336] <= 1'h0;
      write_done_data_log_force[5337] <= 1'h0;
      write_done_data_log_force[5338] <= 1'h0;
      write_done_data_log_force[5339] <= 1'h0;
      write_done_data_log_force[5340] <= 1'h0;
      write_done_data_log_force[5341] <= 1'h0;
      write_done_data_log_force[5342] <= 1'h0;
      write_done_data_log_force[5343] <= 1'h0;
      write_done_data_log_force[5344] <= 1'h0;
      write_done_data_log_force[5345] <= 1'h0;
      write_done_data_log_force[5346] <= 1'h0;
      write_done_data_log_force[5347] <= 1'h0;
      write_done_data_log_force[5348] <= 1'h0;
      write_done_data_log_force[5349] <= 1'h0;
      write_done_data_log_force[5350] <= 1'h0;
      write_done_data_log_force[5351] <= 1'h0;
      write_done_data_log_force[5352] <= 1'h0;
      write_done_data_log_force[5353] <= 1'h0;
      write_done_data_log_force[5354] <= 1'h0;
      write_done_data_log_force[5355] <= 1'h0;
      write_done_data_log_force[5356] <= 1'h0;
      write_done_data_log_force[5357] <= 1'h0;
      write_done_data_log_force[5358] <= 1'h0;
      write_done_data_log_force[5359] <= 1'h0;
      write_done_data_log_force[5360] <= 1'h0;
      write_done_data_log_force[5361] <= 1'h0;
      write_done_data_log_force[5362] <= 1'h0;
      write_done_data_log_force[5363] <= 1'h0;
      write_done_data_log_force[5364] <= 1'h0;
      write_done_data_log_force[5365] <= 1'h0;
      write_done_data_log_force[5366] <= 1'h0;
      write_done_data_log_force[5367] <= 1'h0;
      write_done_data_log_force[5368] <= 1'h0;
      write_done_data_log_force[5369] <= 1'h0;
      write_done_data_log_force[5370] <= 1'h0;
      write_done_data_log_force[5371] <= 1'h0;
      write_done_data_log_force[5372] <= 1'h0;
      write_done_data_log_force[5373] <= 1'h0;
      write_done_data_log_force[5374] <= 1'h0;
      write_done_data_log_force[5375] <= 1'h0;
      write_done_data_log_force[5376] <= 1'h0;
      write_done_data_log_force[5377] <= 1'h0;
      write_done_data_log_force[5378] <= 1'h0;
      write_done_data_log_force[5379] <= 1'h0;
      write_done_data_log_force[5380] <= 1'h0;
      write_done_data_log_force[5381] <= 1'h0;
      write_done_data_log_force[5382] <= 1'h0;
      write_done_data_log_force[5383] <= 1'h0;
      write_done_data_log_force[5384] <= 1'h0;
      write_done_data_log_force[5385] <= 1'h0;
      write_done_data_log_force[5386] <= 1'h0;
      write_done_data_log_force[5387] <= 1'h0;
      write_done_data_log_force[5388] <= 1'h0;
      write_done_data_log_force[5389] <= 1'h0;
      write_done_data_log_force[5390] <= 1'h0;
      write_done_data_log_force[5391] <= 1'h0;
      write_done_data_log_force[5392] <= 1'h0;
      write_done_data_log_force[5393] <= 1'h0;
      write_done_data_log_force[5394] <= 1'h0;
      write_done_data_log_force[5395] <= 1'h0;
      write_done_data_log_force[5396] <= 1'h0;
      write_done_data_log_force[5397] <= 1'h0;
      write_done_data_log_force[5398] <= 1'h0;
      write_done_data_log_force[5399] <= 1'h0;
      write_done_data_log_force[5400] <= 1'h0;
      write_done_data_log_force[5401] <= 1'h0;
      write_done_data_log_force[5402] <= 1'h0;
      write_done_data_log_force[5403] <= 1'h0;
      write_done_data_log_force[5404] <= 1'h0;
      write_done_data_log_force[5405] <= 1'h0;
      write_done_data_log_force[5406] <= 1'h0;
      write_done_data_log_force[5407] <= 1'h0;
      write_done_data_log_force[5408] <= 1'h0;
      write_done_data_log_force[5409] <= 1'h0;
      write_done_data_log_force[5410] <= 1'h0;
      write_done_data_log_force[5411] <= 1'h0;
      write_done_data_log_force[5412] <= 1'h0;
      write_done_data_log_force[5413] <= 1'h0;
      write_done_data_log_force[5414] <= 1'h0;
      write_done_data_log_force[5415] <= 1'h0;
      write_done_data_log_force[5416] <= 1'h0;
      write_done_data_log_force[5417] <= 1'h0;
      write_done_data_log_force[5418] <= 1'h0;
      write_done_data_log_force[5419] <= 1'h0;
      write_done_data_log_force[5420] <= 1'h0;
      write_done_data_log_force[5421] <= 1'h0;
      write_done_data_log_force[5422] <= 1'h0;
      write_done_data_log_force[5423] <= 1'h0;
      write_done_data_log_force[5424] <= 1'h0;
      write_done_data_log_force[5425] <= 1'h0;
      write_done_data_log_force[5426] <= 1'h0;
      write_done_data_log_force[5427] <= 1'h0;
      write_done_data_log_force[5428] <= 1'h0;
      write_done_data_log_force[5429] <= 1'h0;
      write_done_data_log_force[5430] <= 1'h0;
      write_done_data_log_force[5431] <= 1'h0;
      write_done_data_log_force[5432] <= 1'h0;
      write_done_data_log_force[5433] <= 1'h0;
      write_done_data_log_force[5434] <= 1'h0;
      write_done_data_log_force[5435] <= 1'h0;
      write_done_data_log_force[5436] <= 1'h0;
      write_done_data_log_force[5437] <= 1'h0;
      write_done_data_log_force[5438] <= 1'h0;
      write_done_data_log_force[5439] <= 1'h0;
      write_done_data_log_force[5440] <= 1'h0;
      write_done_data_log_force[5441] <= 1'h0;
      write_done_data_log_force[5442] <= 1'h0;
      write_done_data_log_force[5443] <= 1'h0;
      write_done_data_log_force[5444] <= 1'h0;
      write_done_data_log_force[5445] <= 1'h0;
      write_done_data_log_force[5446] <= 1'h0;
      write_done_data_log_force[5447] <= 1'h0;
      write_done_data_log_force[5448] <= 1'h0;
      write_done_data_log_force[5449] <= 1'h0;
      write_done_data_log_force[5450] <= 1'h0;
      write_done_data_log_force[5451] <= 1'h0;
      write_done_data_log_force[5452] <= 1'h0;
      write_done_data_log_force[5453] <= 1'h0;
      write_done_data_log_force[5454] <= 1'h0;
      write_done_data_log_force[5455] <= 1'h0;
      write_done_data_log_force[5456] <= 1'h0;
      write_done_data_log_force[5457] <= 1'h0;
      write_done_data_log_force[5458] <= 1'h0;
      write_done_data_log_force[5459] <= 1'h0;
      write_done_data_log_force[5460] <= 1'h0;
      write_done_data_log_force[5461] <= 1'h0;
      write_done_data_log_force[5462] <= 1'h0;
      write_done_data_log_force[5463] <= 1'h0;
      write_done_data_log_force[5464] <= 1'h0;
      write_done_data_log_force[5465] <= 1'h0;
      write_done_data_log_force[5466] <= 1'h0;
      write_done_data_log_force[5467] <= 1'h0;
      write_done_data_log_force[5468] <= 1'h0;
      write_done_data_log_force[5469] <= 1'h0;
      write_done_data_log_force[5470] <= 1'h0;
      write_done_data_log_force[5471] <= 1'h0;
      write_done_data_log_force[5472] <= 1'h0;
      write_done_data_log_force[5473] <= 1'h0;
      write_done_data_log_force[5474] <= 1'h0;
      write_done_data_log_force[5475] <= 1'h0;
      write_done_data_log_force[5476] <= 1'h0;
      write_done_data_log_force[5477] <= 1'h0;
      write_done_data_log_force[5478] <= 1'h0;
      write_done_data_log_force[5479] <= 1'h0;
      write_done_data_log_force[5480] <= 1'h0;
      write_done_data_log_force[5481] <= 1'h0;
      write_done_data_log_force[5482] <= 1'h0;
      write_done_data_log_force[5483] <= 1'h0;
      write_done_data_log_force[5484] <= 1'h0;
      write_done_data_log_force[5485] <= 1'h0;
      write_done_data_log_force[5486] <= 1'h0;
      write_done_data_log_force[5487] <= 1'h0;
      write_done_data_log_force[5488] <= 1'h0;
      write_done_data_log_force[5489] <= 1'h0;
      write_done_data_log_force[5490] <= 1'h0;
      write_done_data_log_force[5491] <= 1'h0;
      write_done_data_log_force[5492] <= 1'h0;
      write_done_data_log_force[5493] <= 1'h0;
      write_done_data_log_force[5494] <= 1'h0;
      write_done_data_log_force[5495] <= 1'h0;
      write_done_data_log_force[5496] <= 1'h0;
      write_done_data_log_force[5497] <= 1'h0;
      write_done_data_log_force[5498] <= 1'h0;
      write_done_data_log_force[5499] <= 1'h0;
      write_done_data_log_force[5500] <= 1'h0;
      write_done_data_log_force[5501] <= 1'h0;
      write_done_data_log_force[5502] <= 1'h0;
      write_done_data_log_force[5503] <= 1'h0;
      write_done_data_log_force[5504] <= 1'h0;
      write_done_data_log_force[5505] <= 1'h0;
      write_done_data_log_force[5506] <= 1'h0;
      write_done_data_log_force[5507] <= 1'h0;
      write_done_data_log_force[5508] <= 1'h0;
      write_done_data_log_force[5509] <= 1'h0;
      write_done_data_log_force[5510] <= 1'h0;
      write_done_data_log_force[5511] <= 1'h0;
      write_done_data_log_force[5512] <= 1'h0;
      write_done_data_log_force[5513] <= 1'h0;
      write_done_data_log_force[5514] <= 1'h0;
      write_done_data_log_force[5515] <= 1'h0;
      write_done_data_log_force[5516] <= 1'h0;
      write_done_data_log_force[5517] <= 1'h0;
      write_done_data_log_force[5518] <= 1'h0;
      write_done_data_log_force[5519] <= 1'h0;
      write_done_data_log_force[5520] <= 1'h0;
      write_done_data_log_force[5521] <= 1'h0;
      write_done_data_log_force[5522] <= 1'h0;
      write_done_data_log_force[5523] <= 1'h0;
      write_done_data_log_force[5524] <= 1'h0;
      write_done_data_log_force[5525] <= 1'h0;
      write_done_data_log_force[5526] <= 1'h0;
      write_done_data_log_force[5527] <= 1'h0;
      write_done_data_log_force[5528] <= 1'h0;
      write_done_data_log_force[5529] <= 1'h0;
      write_done_data_log_force[5530] <= 1'h0;
      write_done_data_log_force[5531] <= 1'h0;
      write_done_data_log_force[5532] <= 1'h0;
      write_done_data_log_force[5533] <= 1'h0;
      write_done_data_log_force[5534] <= 1'h0;
      write_done_data_log_force[5535] <= 1'h0;
      write_done_data_log_force[5536] <= 1'h0;
      write_done_data_log_force[5537] <= 1'h0;
      write_done_data_log_force[5538] <= 1'h0;
      write_done_data_log_force[5539] <= 1'h0;
      write_done_data_log_force[5540] <= 1'h0;
      write_done_data_log_force[5541] <= 1'h0;
      write_done_data_log_force[5542] <= 1'h0;
      write_done_data_log_force[5543] <= 1'h0;
      write_done_data_log_force[5544] <= 1'h0;
      write_done_data_log_force[5545] <= 1'h0;
      write_done_data_log_force[5546] <= 1'h0;
      write_done_data_log_force[5547] <= 1'h0;
      write_done_data_log_force[5548] <= 1'h0;
      write_done_data_log_force[5549] <= 1'h0;
      write_done_data_log_force[5550] <= 1'h0;
      write_done_data_log_force[5551] <= 1'h0;
      write_done_data_log_force[5552] <= 1'h0;
      write_done_data_log_force[5553] <= 1'h0;
      write_done_data_log_force[5554] <= 1'h0;
      write_done_data_log_force[5555] <= 1'h0;
      write_done_data_log_force[5556] <= 1'h0;
      write_done_data_log_force[5557] <= 1'h0;
      write_done_data_log_force[5558] <= 1'h0;
      write_done_data_log_force[5559] <= 1'h0;
      write_done_data_log_force[5560] <= 1'h0;
      write_done_data_log_force[5561] <= 1'h0;
      write_done_data_log_force[5562] <= 1'h0;
      write_done_data_log_force[5563] <= 1'h0;
      write_done_data_log_force[5564] <= 1'h0;
      write_done_data_log_force[5565] <= 1'h0;
      write_done_data_log_force[5566] <= 1'h0;
      write_done_data_log_force[5567] <= 1'h0;
      write_done_data_log_force[5568] <= 1'h0;
      write_done_data_log_force[5569] <= 1'h0;
      write_done_data_log_force[5570] <= 1'h0;
      write_done_data_log_force[5571] <= 1'h0;
      write_done_data_log_force[5572] <= 1'h0;
      write_done_data_log_force[5573] <= 1'h0;
      write_done_data_log_force[5574] <= 1'h0;
      write_done_data_log_force[5575] <= 1'h0;
      write_done_data_log_force[5576] <= 1'h0;
      write_done_data_log_force[5577] <= 1'h0;
      write_done_data_log_force[5578] <= 1'h0;
      write_done_data_log_force[5579] <= 1'h0;
      write_done_data_log_force[5580] <= 1'h0;
      write_done_data_log_force[5581] <= 1'h0;
      write_done_data_log_force[5582] <= 1'h0;
      write_done_data_log_force[5583] <= 1'h0;
      write_done_data_log_force[5584] <= 1'h0;
      write_done_data_log_force[5585] <= 1'h0;
      write_done_data_log_force[5586] <= 1'h0;
      write_done_data_log_force[5587] <= 1'h0;
      write_done_data_log_force[5588] <= 1'h0;
      write_done_data_log_force[5589] <= 1'h0;
      write_done_data_log_force[5590] <= 1'h0;
      write_done_data_log_force[5591] <= 1'h0;
      write_done_data_log_force[5592] <= 1'h0;
      write_done_data_log_force[5593] <= 1'h0;
      write_done_data_log_force[5594] <= 1'h0;
      write_done_data_log_force[5595] <= 1'h0;
      write_done_data_log_force[5596] <= 1'h0;
      write_done_data_log_force[5597] <= 1'h0;
      write_done_data_log_force[5598] <= 1'h0;
      write_done_data_log_force[5599] <= 1'h0;
      write_done_data_log_force[5600] <= 1'h0;
      write_done_data_log_force[5601] <= 1'h0;
      write_done_data_log_force[5602] <= 1'h0;
      write_done_data_log_force[5603] <= 1'h0;
      write_done_data_log_force[5604] <= 1'h0;
      write_done_data_log_force[5605] <= 1'h0;
      write_done_data_log_force[5606] <= 1'h0;
      write_done_data_log_force[5607] <= 1'h0;
      write_done_data_log_force[5608] <= 1'h0;
      write_done_data_log_force[5609] <= 1'h0;
      write_done_data_log_force[5610] <= 1'h0;
      write_done_data_log_force[5611] <= 1'h0;
      write_done_data_log_force[5612] <= 1'h0;
      write_done_data_log_force[5613] <= 1'h0;
      write_done_data_log_force[5614] <= 1'h0;
      write_done_data_log_force[5615] <= 1'h0;
      write_done_data_log_force[5616] <= 1'h0;
      write_done_data_log_force[5617] <= 1'h0;
      write_done_data_log_force[5618] <= 1'h0;
      write_done_data_log_force[5619] <= 1'h0;
      write_done_data_log_force[5620] <= 1'h0;
      write_done_data_log_force[5621] <= 1'h0;
      write_done_data_log_force[5622] <= 1'h0;
      write_done_data_log_force[5623] <= 1'h0;
      write_done_data_log_force[5624] <= 1'h0;
      write_done_data_log_force[5625] <= 1'h0;
      write_done_data_log_force[5626] <= 1'h0;
      write_done_data_log_force[5627] <= 1'h0;
      write_done_data_log_force[5628] <= 1'h0;
      write_done_data_log_force[5629] <= 1'h0;
      write_done_data_log_force[5630] <= 1'h0;
      write_done_data_log_force[5631] <= 1'h0;
      write_done_data_log_force[5632] <= 1'h0;
      write_done_data_log_force[5633] <= 1'h0;
      write_done_data_log_force[5634] <= 1'h0;
      write_done_data_log_force[5635] <= 1'h0;
      write_done_data_log_force[5636] <= 1'h0;
      write_done_data_log_force[5637] <= 1'h0;
      write_done_data_log_force[5638] <= 1'h0;
      write_done_data_log_force[5639] <= 1'h0;
      write_done_data_log_force[5640] <= 1'h0;
      write_done_data_log_force[5641] <= 1'h0;
      write_done_data_log_force[5642] <= 1'h0;
      write_done_data_log_force[5643] <= 1'h0;
      write_done_data_log_force[5644] <= 1'h0;
      write_done_data_log_force[5645] <= 1'h0;
      write_done_data_log_force[5646] <= 1'h0;
      write_done_data_log_force[5647] <= 1'h0;
      write_done_data_log_force[5648] <= 1'h0;
      write_done_data_log_force[5649] <= 1'h0;
      write_done_data_log_force[5650] <= 1'h0;
      write_done_data_log_force[5651] <= 1'h0;
      write_done_data_log_force[5652] <= 1'h0;
      write_done_data_log_force[5653] <= 1'h0;
      write_done_data_log_force[5654] <= 1'h0;
      write_done_data_log_force[5655] <= 1'h0;
      write_done_data_log_force[5656] <= 1'h0;
      write_done_data_log_force[5657] <= 1'h0;
      write_done_data_log_force[5658] <= 1'h0;
      write_done_data_log_force[5659] <= 1'h0;
      write_done_data_log_force[5660] <= 1'h0;
      write_done_data_log_force[5661] <= 1'h0;
      write_done_data_log_force[5662] <= 1'h0;
      write_done_data_log_force[5663] <= 1'h0;
      write_done_data_log_force[5664] <= 1'h0;
      write_done_data_log_force[5665] <= 1'h0;
      write_done_data_log_force[5666] <= 1'h0;
      write_done_data_log_force[5667] <= 1'h0;
      write_done_data_log_force[5668] <= 1'h0;
      write_done_data_log_force[5669] <= 1'h0;
      write_done_data_log_force[5670] <= 1'h0;
      write_done_data_log_force[5671] <= 1'h0;
      write_done_data_log_force[5672] <= 1'h0;
      write_done_data_log_force[5673] <= 1'h0;
      write_done_data_log_force[5674] <= 1'h0;
      write_done_data_log_force[5675] <= 1'h0;
      write_done_data_log_force[5676] <= 1'h0;
      write_done_data_log_force[5677] <= 1'h0;
      write_done_data_log_force[5678] <= 1'h0;
      write_done_data_log_force[5679] <= 1'h0;
      write_done_data_log_force[5680] <= 1'h0;
      write_done_data_log_force[5681] <= 1'h0;
      write_done_data_log_force[5682] <= 1'h0;
      write_done_data_log_force[5683] <= 1'h0;
      write_done_data_log_force[5684] <= 1'h0;
      write_done_data_log_force[5685] <= 1'h0;
      write_done_data_log_force[5686] <= 1'h0;
      write_done_data_log_force[5687] <= 1'h0;
      write_done_data_log_force[5688] <= 1'h0;
      write_done_data_log_force[5689] <= 1'h0;
      write_done_data_log_force[5690] <= 1'h0;
      write_done_data_log_force[5691] <= 1'h0;
      write_done_data_log_force[5692] <= 1'h0;
      write_done_data_log_force[5693] <= 1'h0;
      write_done_data_log_force[5694] <= 1'h0;
      write_done_data_log_force[5695] <= 1'h0;
      write_done_data_log_force[5696] <= 1'h0;
      write_done_data_log_force[5697] <= 1'h0;
      write_done_data_log_force[5698] <= 1'h0;
      write_done_data_log_force[5699] <= 1'h0;
      write_done_data_log_force[5700] <= 1'h0;
      write_done_data_log_force[5701] <= 1'h0;
      write_done_data_log_force[5702] <= 1'h0;
      write_done_data_log_force[5703] <= 1'h0;
      write_done_data_log_force[5704] <= 1'h0;
      write_done_data_log_force[5705] <= 1'h0;
      write_done_data_log_force[5706] <= 1'h0;
      write_done_data_log_force[5707] <= 1'h0;
      write_done_data_log_force[5708] <= 1'h0;
      write_done_data_log_force[5709] <= 1'h0;
      write_done_data_log_force[5710] <= 1'h0;
      write_done_data_log_force[5711] <= 1'h0;
      write_done_data_log_force[5712] <= 1'h0;
      write_done_data_log_force[5713] <= 1'h0;
      write_done_data_log_force[5714] <= 1'h0;
      write_done_data_log_force[5715] <= 1'h0;
      write_done_data_log_force[5716] <= 1'h0;
      write_done_data_log_force[5717] <= 1'h0;
      write_done_data_log_force[5718] <= 1'h0;
      write_done_data_log_force[5719] <= 1'h0;
      write_done_data_log_force[5720] <= 1'h0;
      write_done_data_log_force[5721] <= 1'h0;
      write_done_data_log_force[5722] <= 1'h0;
      write_done_data_log_force[5723] <= 1'h0;
      write_done_data_log_force[5724] <= 1'h0;
      write_done_data_log_force[5725] <= 1'h0;
      write_done_data_log_force[5726] <= 1'h0;
      write_done_data_log_force[5727] <= 1'h0;
      write_done_data_log_force[5728] <= 1'h0;
      write_done_data_log_force[5729] <= 1'h0;
      write_done_data_log_force[5730] <= 1'h0;
      write_done_data_log_force[5731] <= 1'h0;
      write_done_data_log_force[5732] <= 1'h0;
      write_done_data_log_force[5733] <= 1'h0;
      write_done_data_log_force[5734] <= 1'h0;
      write_done_data_log_force[5735] <= 1'h0;
      write_done_data_log_force[5736] <= 1'h0;
      write_done_data_log_force[5737] <= 1'h0;
      write_done_data_log_force[5738] <= 1'h0;
      write_done_data_log_force[5739] <= 1'h0;
      write_done_data_log_force[5740] <= 1'h0;
      write_done_data_log_force[5741] <= 1'h0;
      write_done_data_log_force[5742] <= 1'h0;
      write_done_data_log_force[5743] <= 1'h0;
      write_done_data_log_force[5744] <= 1'h0;
      write_done_data_log_force[5745] <= 1'h0;
      write_done_data_log_force[5746] <= 1'h0;
      write_done_data_log_force[5747] <= 1'h0;
      write_done_data_log_force[5748] <= 1'h0;
      write_done_data_log_force[5749] <= 1'h0;
      write_done_data_log_force[5750] <= 1'h0;
      write_done_data_log_force[5751] <= 1'h0;
      write_done_data_log_force[5752] <= 1'h0;
      write_done_data_log_force[5753] <= 1'h0;
      write_done_data_log_force[5754] <= 1'h0;
      write_done_data_log_force[5755] <= 1'h0;
      write_done_data_log_force[5756] <= 1'h0;
      write_done_data_log_force[5757] <= 1'h0;
      write_done_data_log_force[5758] <= 1'h0;
      write_done_data_log_force[5759] <= 1'h0;
      write_done_data_log_force[5760] <= 1'h0;
      write_done_data_log_force[5761] <= 1'h0;
      write_done_data_log_force[5762] <= 1'h0;
      write_done_data_log_force[5763] <= 1'h0;
      write_done_data_log_force[5764] <= 1'h0;
      write_done_data_log_force[5765] <= 1'h0;
      write_done_data_log_force[5766] <= 1'h0;
      write_done_data_log_force[5767] <= 1'h0;
      write_done_data_log_force[5768] <= 1'h0;
      write_done_data_log_force[5769] <= 1'h0;
      write_done_data_log_force[5770] <= 1'h0;
      write_done_data_log_force[5771] <= 1'h0;
      write_done_data_log_force[5772] <= 1'h0;
      write_done_data_log_force[5773] <= 1'h0;
      write_done_data_log_force[5774] <= 1'h0;
      write_done_data_log_force[5775] <= 1'h0;
      write_done_data_log_force[5776] <= 1'h0;
      write_done_data_log_force[5777] <= 1'h0;
      write_done_data_log_force[5778] <= 1'h0;
      write_done_data_log_force[5779] <= 1'h0;
      write_done_data_log_force[5780] <= 1'h0;
      write_done_data_log_force[5781] <= 1'h0;
      write_done_data_log_force[5782] <= 1'h0;
      write_done_data_log_force[5783] <= 1'h0;
      write_done_data_log_force[5784] <= 1'h0;
      write_done_data_log_force[5785] <= 1'h0;
      write_done_data_log_force[5786] <= 1'h0;
      write_done_data_log_force[5787] <= 1'h0;
      write_done_data_log_force[5788] <= 1'h0;
      write_done_data_log_force[5789] <= 1'h0;
      write_done_data_log_force[5790] <= 1'h0;
      write_done_data_log_force[5791] <= 1'h0;
      write_done_data_log_force[5792] <= 1'h0;
      write_done_data_log_force[5793] <= 1'h0;
      write_done_data_log_force[5794] <= 1'h0;
      write_done_data_log_force[5795] <= 1'h0;
      write_done_data_log_force[5796] <= 1'h0;
      write_done_data_log_force[5797] <= 1'h0;
      write_done_data_log_force[5798] <= 1'h0;
      write_done_data_log_force[5799] <= 1'h0;
      write_done_data_log_force[5800] <= 1'h0;
      write_done_data_log_force[5801] <= 1'h0;
      write_done_data_log_force[5802] <= 1'h0;
      write_done_data_log_force[5803] <= 1'h0;
      write_done_data_log_force[5804] <= 1'h0;
      write_done_data_log_force[5805] <= 1'h0;
      write_done_data_log_force[5806] <= 1'h0;
      write_done_data_log_force[5807] <= 1'h0;
      write_done_data_log_force[5808] <= 1'h0;
      write_done_data_log_force[5809] <= 1'h0;
      write_done_data_log_force[5810] <= 1'h0;
      write_done_data_log_force[5811] <= 1'h0;
      write_done_data_log_force[5812] <= 1'h0;
      write_done_data_log_force[5813] <= 1'h0;
      write_done_data_log_force[5814] <= 1'h0;
      write_done_data_log_force[5815] <= 1'h0;
      write_done_data_log_force[5816] <= 1'h0;
      write_done_data_log_force[5817] <= 1'h0;
      write_done_data_log_force[5818] <= 1'h0;
      write_done_data_log_force[5819] <= 1'h0;
      write_done_data_log_force[5820] <= 1'h0;
      write_done_data_log_force[5821] <= 1'h0;
      write_done_data_log_force[5822] <= 1'h0;
      write_done_data_log_force[5823] <= 1'h0;
      write_done_data_log_force[5824] <= 1'h0;
      write_done_data_log_force[5825] <= 1'h0;
      write_done_data_log_force[5826] <= 1'h0;
      write_done_data_log_force[5827] <= 1'h0;
      write_done_data_log_force[5828] <= 1'h0;
      write_done_data_log_force[5829] <= 1'h0;
      write_done_data_log_force[5830] <= 1'h0;
      write_done_data_log_force[5831] <= 1'h0;
      write_done_data_log_force[5832] <= 1'h0;
      write_done_data_log_force[5833] <= 1'h0;
      write_done_data_log_force[5834] <= 1'h0;
      write_done_data_log_force[5835] <= 1'h0;
      write_done_data_log_force[5836] <= 1'h0;
      write_done_data_log_force[5837] <= 1'h0;
      write_done_data_log_force[5838] <= 1'h0;
      write_done_data_log_force[5839] <= 1'h0;
      write_done_data_log_force[5840] <= 1'h0;
      write_done_data_log_force[5841] <= 1'h0;
      write_done_data_log_force[5842] <= 1'h0;
      write_done_data_log_force[5843] <= 1'h0;
      write_done_data_log_force[5844] <= 1'h0;
      write_done_data_log_force[5845] <= 1'h0;
      write_done_data_log_force[5846] <= 1'h0;
      write_done_data_log_force[5847] <= 1'h0;
      write_done_data_log_force[5848] <= 1'h0;
      write_done_data_log_force[5849] <= 1'h0;
      write_done_data_log_force[5850] <= 1'h0;
      write_done_data_log_force[5851] <= 1'h0;
      write_done_data_log_force[5852] <= 1'h0;
      write_done_data_log_force[5853] <= 1'h0;
      write_done_data_log_force[5854] <= 1'h0;
      write_done_data_log_force[5855] <= 1'h0;
      write_done_data_log_force[5856] <= 1'h0;
      write_done_data_log_force[5857] <= 1'h0;
      write_done_data_log_force[5858] <= 1'h0;
      write_done_data_log_force[5859] <= 1'h0;
      write_done_data_log_force[5860] <= 1'h0;
      write_done_data_log_force[5861] <= 1'h0;
      write_done_data_log_force[5862] <= 1'h0;
      write_done_data_log_force[5863] <= 1'h0;
      write_done_data_log_force[5864] <= 1'h0;
      write_done_data_log_force[5865] <= 1'h0;
      write_done_data_log_force[5866] <= 1'h0;
      write_done_data_log_force[5867] <= 1'h0;
      write_done_data_log_force[5868] <= 1'h0;
      write_done_data_log_force[5869] <= 1'h0;
      write_done_data_log_force[5870] <= 1'h0;
      write_done_data_log_force[5871] <= 1'h0;
      write_done_data_log_force[5872] <= 1'h0;
      write_done_data_log_force[5873] <= 1'h0;
      write_done_data_log_force[5874] <= 1'h0;
      write_done_data_log_force[5875] <= 1'h0;
      write_done_data_log_force[5876] <= 1'h0;
      write_done_data_log_force[5877] <= 1'h0;
      write_done_data_log_force[5878] <= 1'h0;
      write_done_data_log_force[5879] <= 1'h0;
      write_done_data_log_force[5880] <= 1'h0;
      write_done_data_log_force[5881] <= 1'h0;
      write_done_data_log_force[5882] <= 1'h0;
      write_done_data_log_force[5883] <= 1'h0;
      write_done_data_log_force[5884] <= 1'h0;
      write_done_data_log_force[5885] <= 1'h0;
      write_done_data_log_force[5886] <= 1'h0;
      write_done_data_log_force[5887] <= 1'h0;
      write_done_data_log_force[5888] <= 1'h0;
      write_done_data_log_force[5889] <= 1'h0;
      write_done_data_log_force[5890] <= 1'h0;
      write_done_data_log_force[5891] <= 1'h0;
      write_done_data_log_force[5892] <= 1'h0;
      write_done_data_log_force[5893] <= 1'h0;
      write_done_data_log_force[5894] <= 1'h0;
      write_done_data_log_force[5895] <= 1'h0;
      write_done_data_log_force[5896] <= 1'h0;
      write_done_data_log_force[5897] <= 1'h0;
      write_done_data_log_force[5898] <= 1'h0;
      write_done_data_log_force[5899] <= 1'h0;
      write_done_data_log_force[5900] <= 1'h0;
      write_done_data_log_force[5901] <= 1'h0;
      write_done_data_log_force[5902] <= 1'h0;
      write_done_data_log_force[5903] <= 1'h0;
      write_done_data_log_force[5904] <= 1'h0;
      write_done_data_log_force[5905] <= 1'h0;
      write_done_data_log_force[5906] <= 1'h0;
      write_done_data_log_force[5907] <= 1'h0;
      write_done_data_log_force[5908] <= 1'h0;
      write_done_data_log_force[5909] <= 1'h0;
      write_done_data_log_force[5910] <= 1'h0;
      write_done_data_log_force[5911] <= 1'h0;
      write_done_data_log_force[5912] <= 1'h0;
      write_done_data_log_force[5913] <= 1'h0;
      write_done_data_log_force[5914] <= 1'h0;
      write_done_data_log_force[5915] <= 1'h0;
      write_done_data_log_force[5916] <= 1'h0;
      write_done_data_log_force[5917] <= 1'h0;
      write_done_data_log_force[5918] <= 1'h0;
      write_done_data_log_force[5919] <= 1'h0;
      write_done_data_log_force[5920] <= 1'h0;
      write_done_data_log_force[5921] <= 1'h0;
      write_done_data_log_force[5922] <= 1'h0;
      write_done_data_log_force[5923] <= 1'h0;
      write_done_data_log_force[5924] <= 1'h0;
      write_done_data_log_force[5925] <= 1'h0;
      write_done_data_log_force[5926] <= 1'h0;
      write_done_data_log_force[5927] <= 1'h0;
      write_done_data_log_force[5928] <= 1'h0;
      write_done_data_log_force[5929] <= 1'h0;
      write_done_data_log_force[5930] <= 1'h0;
      write_done_data_log_force[5931] <= 1'h0;
      write_done_data_log_force[5932] <= 1'h0;
      write_done_data_log_force[5933] <= 1'h0;
      write_done_data_log_force[5934] <= 1'h0;
      write_done_data_log_force[5935] <= 1'h0;
      write_done_data_log_force[5936] <= 1'h0;
      write_done_data_log_force[5937] <= 1'h0;
      write_done_data_log_force[5938] <= 1'h0;
      write_done_data_log_force[5939] <= 1'h0;
      write_done_data_log_force[5940] <= 1'h0;
      write_done_data_log_force[5941] <= 1'h0;
      write_done_data_log_force[5942] <= 1'h0;
      write_done_data_log_force[5943] <= 1'h0;
      write_done_data_log_force[5944] <= 1'h0;
      write_done_data_log_force[5945] <= 1'h0;
      write_done_data_log_force[5946] <= 1'h0;
      write_done_data_log_force[5947] <= 1'h0;
      write_done_data_log_force[5948] <= 1'h0;
      write_done_data_log_force[5949] <= 1'h0;
      write_done_data_log_force[5950] <= 1'h0;
      write_done_data_log_force[5951] <= 1'h0;
      write_done_data_log_force[5952] <= 1'h0;
      write_done_data_log_force[5953] <= 1'h0;
      write_done_data_log_force[5954] <= 1'h0;
      write_done_data_log_force[5955] <= 1'h0;
      write_done_data_log_force[5956] <= 1'h0;
      write_done_data_log_force[5957] <= 1'h0;
      write_done_data_log_force[5958] <= 1'h0;
      write_done_data_log_force[5959] <= 1'h0;
      write_done_data_log_force[5960] <= 1'h0;
      write_done_data_log_force[5961] <= 1'h0;
      write_done_data_log_force[5962] <= 1'h0;
      write_done_data_log_force[5963] <= 1'h0;
      write_done_data_log_force[5964] <= 1'h0;
      write_done_data_log_force[5965] <= 1'h0;
      write_done_data_log_force[5966] <= 1'h0;
      write_done_data_log_force[5967] <= 1'h0;
      write_done_data_log_force[5968] <= 1'h0;
      write_done_data_log_force[5969] <= 1'h0;
      write_done_data_log_force[5970] <= 1'h0;
      write_done_data_log_force[5971] <= 1'h0;
      write_done_data_log_force[5972] <= 1'h0;
      write_done_data_log_force[5973] <= 1'h0;
      write_done_data_log_force[5974] <= 1'h0;
      write_done_data_log_force[5975] <= 1'h0;
      write_done_data_log_force[5976] <= 1'h0;
      write_done_data_log_force[5977] <= 1'h0;
      write_done_data_log_force[5978] <= 1'h0;
      write_done_data_log_force[5979] <= 1'h0;
      write_done_data_log_force[5980] <= 1'h0;
      write_done_data_log_force[5981] <= 1'h0;
      write_done_data_log_force[5982] <= 1'h0;
      write_done_data_log_force[5983] <= 1'h0;
      write_done_data_log_force[5984] <= 1'h0;
      write_done_data_log_force[5985] <= 1'h0;
      write_done_data_log_force[5986] <= 1'h0;
      write_done_data_log_force[5987] <= 1'h0;
      write_done_data_log_force[5988] <= 1'h0;
      write_done_data_log_force[5989] <= 1'h0;
      write_done_data_log_force[5990] <= 1'h0;
      write_done_data_log_force[5991] <= 1'h0;
      write_done_data_log_force[5992] <= 1'h0;
      write_done_data_log_force[5993] <= 1'h0;
      write_done_data_log_force[5994] <= 1'h0;
      write_done_data_log_force[5995] <= 1'h0;
      write_done_data_log_force[5996] <= 1'h0;
      write_done_data_log_force[5997] <= 1'h0;
      write_done_data_log_force[5998] <= 1'h0;
      write_done_data_log_force[5999] <= 1'h0;
      write_done_data_log_force[6000] <= 1'h0;
      write_done_data_log_force[6001] <= 1'h0;
      write_done_data_log_force[6002] <= 1'h0;
      write_done_data_log_force[6003] <= 1'h0;
      write_done_data_log_force[6004] <= 1'h0;
      write_done_data_log_force[6005] <= 1'h0;
      write_done_data_log_force[6006] <= 1'h0;
      write_done_data_log_force[6007] <= 1'h0;
      write_done_data_log_force[6008] <= 1'h0;
      write_done_data_log_force[6009] <= 1'h0;
      write_done_data_log_force[6010] <= 1'h0;
      write_done_data_log_force[6011] <= 1'h0;
      write_done_data_log_force[6012] <= 1'h0;
      write_done_data_log_force[6013] <= 1'h0;
      write_done_data_log_force[6014] <= 1'h0;
      write_done_data_log_force[6015] <= 1'h0;
      write_done_data_log_force[6016] <= 1'h0;
      write_done_data_log_force[6017] <= 1'h0;
      write_done_data_log_force[6018] <= 1'h0;
      write_done_data_log_force[6019] <= 1'h0;
      write_done_data_log_force[6020] <= 1'h0;
      write_done_data_log_force[6021] <= 1'h0;
      write_done_data_log_force[6022] <= 1'h0;
      write_done_data_log_force[6023] <= 1'h0;
      write_done_data_log_force[6024] <= 1'h0;
      write_done_data_log_force[6025] <= 1'h0;
      write_done_data_log_force[6026] <= 1'h0;
      write_done_data_log_force[6027] <= 1'h0;
      write_done_data_log_force[6028] <= 1'h0;
      write_done_data_log_force[6029] <= 1'h0;
      write_done_data_log_force[6030] <= 1'h0;
      write_done_data_log_force[6031] <= 1'h0;
      write_done_data_log_force[6032] <= 1'h0;
      write_done_data_log_force[6033] <= 1'h0;
      write_done_data_log_force[6034] <= 1'h0;
      write_done_data_log_force[6035] <= 1'h0;
      write_done_data_log_force[6036] <= 1'h0;
      write_done_data_log_force[6037] <= 1'h0;
      write_done_data_log_force[6038] <= 1'h0;
      write_done_data_log_force[6039] <= 1'h0;
      write_done_data_log_force[6040] <= 1'h0;
      write_done_data_log_force[6041] <= 1'h0;
      write_done_data_log_force[6042] <= 1'h0;
      write_done_data_log_force[6043] <= 1'h0;
      write_done_data_log_force[6044] <= 1'h0;
      write_done_data_log_force[6045] <= 1'h0;
      write_done_data_log_force[6046] <= 1'h0;
      write_done_data_log_force[6047] <= 1'h0;
      write_done_data_log_force[6048] <= 1'h0;
      write_done_data_log_force[6049] <= 1'h0;
      write_done_data_log_force[6050] <= 1'h0;
      write_done_data_log_force[6051] <= 1'h0;
      write_done_data_log_force[6052] <= 1'h0;
      write_done_data_log_force[6053] <= 1'h0;
      write_done_data_log_force[6054] <= 1'h0;
      write_done_data_log_force[6055] <= 1'h0;
      write_done_data_log_force[6056] <= 1'h0;
      write_done_data_log_force[6057] <= 1'h0;
      write_done_data_log_force[6058] <= 1'h0;
      write_done_data_log_force[6059] <= 1'h0;
      write_done_data_log_force[6060] <= 1'h0;
      write_done_data_log_force[6061] <= 1'h0;
      write_done_data_log_force[6062] <= 1'h0;
      write_done_data_log_force[6063] <= 1'h0;
      write_done_data_log_force[6064] <= 1'h0;
      write_done_data_log_force[6065] <= 1'h0;
      write_done_data_log_force[6066] <= 1'h0;
      write_done_data_log_force[6067] <= 1'h0;
      write_done_data_log_force[6068] <= 1'h0;
      write_done_data_log_force[6069] <= 1'h0;
      write_done_data_log_force[6070] <= 1'h0;
      write_done_data_log_force[6071] <= 1'h0;
      write_done_data_log_force[6072] <= 1'h0;
      write_done_data_log_force[6073] <= 1'h0;
      write_done_data_log_force[6074] <= 1'h0;
      write_done_data_log_force[6075] <= 1'h0;
      write_done_data_log_force[6076] <= 1'h0;
      write_done_data_log_force[6077] <= 1'h0;
      write_done_data_log_force[6078] <= 1'h0;
      write_done_data_log_force[6079] <= 1'h0;
      write_done_data_log_force[6080] <= 1'h0;
      write_done_data_log_force[6081] <= 1'h0;
      write_done_data_log_force[6082] <= 1'h0;
      write_done_data_log_force[6083] <= 1'h0;
      write_done_data_log_force[6084] <= 1'h0;
      write_done_data_log_force[6085] <= 1'h0;
      write_done_data_log_force[6086] <= 1'h0;
      write_done_data_log_force[6087] <= 1'h0;
      write_done_data_log_force[6088] <= 1'h0;
      write_done_data_log_force[6089] <= 1'h0;
      write_done_data_log_force[6090] <= 1'h0;
      write_done_data_log_force[6091] <= 1'h0;
      write_done_data_log_force[6092] <= 1'h0;
      write_done_data_log_force[6093] <= 1'h0;
      write_done_data_log_force[6094] <= 1'h0;
      write_done_data_log_force[6095] <= 1'h0;
      write_done_data_log_force[6096] <= 1'h0;
      write_done_data_log_force[6097] <= 1'h0;
      write_done_data_log_force[6098] <= 1'h0;
      write_done_data_log_force[6099] <= 1'h0;
      write_done_data_log_force[6100] <= 1'h0;
      write_done_data_log_force[6101] <= 1'h0;
      write_done_data_log_force[6102] <= 1'h0;
      write_done_data_log_force[6103] <= 1'h0;
      write_done_data_log_force[6104] <= 1'h0;
      write_done_data_log_force[6105] <= 1'h0;
      write_done_data_log_force[6106] <= 1'h0;
      write_done_data_log_force[6107] <= 1'h0;
      write_done_data_log_force[6108] <= 1'h0;
      write_done_data_log_force[6109] <= 1'h0;
      write_done_data_log_force[6110] <= 1'h0;
      write_done_data_log_force[6111] <= 1'h0;
      write_done_data_log_force[6112] <= 1'h0;
      write_done_data_log_force[6113] <= 1'h0;
      write_done_data_log_force[6114] <= 1'h0;
      write_done_data_log_force[6115] <= 1'h0;
      write_done_data_log_force[6116] <= 1'h0;
      write_done_data_log_force[6117] <= 1'h0;
      write_done_data_log_force[6118] <= 1'h0;
      write_done_data_log_force[6119] <= 1'h0;
      write_done_data_log_force[6120] <= 1'h0;
      write_done_data_log_force[6121] <= 1'h0;
      write_done_data_log_force[6122] <= 1'h0;
      write_done_data_log_force[6123] <= 1'h0;
      write_done_data_log_force[6124] <= 1'h0;
      write_done_data_log_force[6125] <= 1'h0;
      write_done_data_log_force[6126] <= 1'h0;
      write_done_data_log_force[6127] <= 1'h0;
      write_done_data_log_force[6128] <= 1'h0;
      write_done_data_log_force[6129] <= 1'h0;
      write_done_data_log_force[6130] <= 1'h0;
      write_done_data_log_force[6131] <= 1'h0;
      write_done_data_log_force[6132] <= 1'h0;
      write_done_data_log_force[6133] <= 1'h0;
      write_done_data_log_force[6134] <= 1'h0;
      write_done_data_log_force[6135] <= 1'h0;
      write_done_data_log_force[6136] <= 1'h0;
      write_done_data_log_force[6137] <= 1'h0;
      write_done_data_log_force[6138] <= 1'h0;
      write_done_data_log_force[6139] <= 1'h0;
      write_done_data_log_force[6140] <= 1'h0;
      write_done_data_log_force[6141] <= 1'h0;
      write_done_data_log_force[6142] <= 1'h0;
      write_done_data_log_force[6143] <= 1'h0;
      write_done_data_log_force[6144] <= 1'h0;
      write_done_data_log_force[6145] <= 1'h0;
      write_done_data_log_force[6146] <= 1'h0;
      write_done_data_log_force[6147] <= 1'h0;
      write_done_data_log_force[6148] <= 1'h0;
      write_done_data_log_force[6149] <= 1'h0;
      write_done_data_log_force[6150] <= 1'h0;
      write_done_data_log_force[6151] <= 1'h0;
      write_done_data_log_force[6152] <= 1'h0;
      write_done_data_log_force[6153] <= 1'h0;
      write_done_data_log_force[6154] <= 1'h0;
      write_done_data_log_force[6155] <= 1'h0;
      write_done_data_log_force[6156] <= 1'h0;
      write_done_data_log_force[6157] <= 1'h0;
      write_done_data_log_force[6158] <= 1'h0;
      write_done_data_log_force[6159] <= 1'h0;
      write_done_data_log_force[6160] <= 1'h0;
      write_done_data_log_force[6161] <= 1'h0;
      write_done_data_log_force[6162] <= 1'h0;
      write_done_data_log_force[6163] <= 1'h0;
      write_done_data_log_force[6164] <= 1'h0;
      write_done_data_log_force[6165] <= 1'h0;
      write_done_data_log_force[6166] <= 1'h0;
      write_done_data_log_force[6167] <= 1'h0;
      write_done_data_log_force[6168] <= 1'h0;
      write_done_data_log_force[6169] <= 1'h0;
      write_done_data_log_force[6170] <= 1'h0;
      write_done_data_log_force[6171] <= 1'h0;
      write_done_data_log_force[6172] <= 1'h0;
      write_done_data_log_force[6173] <= 1'h0;
      write_done_data_log_force[6174] <= 1'h0;
      write_done_data_log_force[6175] <= 1'h0;
      write_done_data_log_force[6176] <= 1'h0;
      write_done_data_log_force[6177] <= 1'h0;
      write_done_data_log_force[6178] <= 1'h0;
      write_done_data_log_force[6179] <= 1'h0;
      write_done_data_log_force[6180] <= 1'h0;
      write_done_data_log_force[6181] <= 1'h0;
      write_done_data_log_force[6182] <= 1'h0;
      write_done_data_log_force[6183] <= 1'h0;
      write_done_data_log_force[6184] <= 1'h0;
      write_done_data_log_force[6185] <= 1'h0;
      write_done_data_log_force[6186] <= 1'h0;
      write_done_data_log_force[6187] <= 1'h0;
      write_done_data_log_force[6188] <= 1'h0;
      write_done_data_log_force[6189] <= 1'h0;
      write_done_data_log_force[6190] <= 1'h0;
      write_done_data_log_force[6191] <= 1'h0;
      write_done_data_log_force[6192] <= 1'h0;
      write_done_data_log_force[6193] <= 1'h0;
      write_done_data_log_force[6194] <= 1'h0;
      write_done_data_log_force[6195] <= 1'h0;
      write_done_data_log_force[6196] <= 1'h0;
      write_done_data_log_force[6197] <= 1'h0;
      write_done_data_log_force[6198] <= 1'h0;
      write_done_data_log_force[6199] <= 1'h0;
      write_done_data_log_force[6200] <= 1'h0;
      write_done_data_log_force[6201] <= 1'h0;
      write_done_data_log_force[6202] <= 1'h0;
      write_done_data_log_force[6203] <= 1'h0;
      write_done_data_log_force[6204] <= 1'h0;
      write_done_data_log_force[6205] <= 1'h0;
      write_done_data_log_force[6206] <= 1'h0;
      write_done_data_log_force[6207] <= 1'h0;
      write_done_data_log_force[6208] <= 1'h0;
      write_done_data_log_force[6209] <= 1'h0;
      write_done_data_log_force[6210] <= 1'h0;
      write_done_data_log_force[6211] <= 1'h0;
      write_done_data_log_force[6212] <= 1'h0;
      write_done_data_log_force[6213] <= 1'h0;
      write_done_data_log_force[6214] <= 1'h0;
      write_done_data_log_force[6215] <= 1'h0;
      write_done_data_log_force[6216] <= 1'h0;
      write_done_data_log_force[6217] <= 1'h0;
      write_done_data_log_force[6218] <= 1'h0;
      write_done_data_log_force[6219] <= 1'h0;
      write_done_data_log_force[6220] <= 1'h0;
      write_done_data_log_force[6221] <= 1'h0;
      write_done_data_log_force[6222] <= 1'h0;
      write_done_data_log_force[6223] <= 1'h0;
      write_done_data_log_force[6224] <= 1'h0;
      write_done_data_log_force[6225] <= 1'h0;
      write_done_data_log_force[6226] <= 1'h0;
      write_done_data_log_force[6227] <= 1'h0;
      write_done_data_log_force[6228] <= 1'h0;
      write_done_data_log_force[6229] <= 1'h0;
      write_done_data_log_force[6230] <= 1'h0;
      write_done_data_log_force[6231] <= 1'h0;
      write_done_data_log_force[6232] <= 1'h0;
      write_done_data_log_force[6233] <= 1'h0;
      write_done_data_log_force[6234] <= 1'h0;
      write_done_data_log_force[6235] <= 1'h0;
      write_done_data_log_force[6236] <= 1'h0;
      write_done_data_log_force[6237] <= 1'h0;
      write_done_data_log_force[6238] <= 1'h0;
      write_done_data_log_force[6239] <= 1'h0;
      write_done_data_log_force[6240] <= 1'h0;
      write_done_data_log_force[6241] <= 1'h0;
      write_done_data_log_force[6242] <= 1'h0;
      write_done_data_log_force[6243] <= 1'h0;
      write_done_data_log_force[6244] <= 1'h0;
      write_done_data_log_force[6245] <= 1'h0;
      write_done_data_log_force[6246] <= 1'h0;
      write_done_data_log_force[6247] <= 1'h0;
      write_done_data_log_force[6248] <= 1'h0;
      write_done_data_log_force[6249] <= 1'h0;
      write_done_data_log_force[6250] <= 1'h0;
      write_done_data_log_force[6251] <= 1'h0;
      write_done_data_log_force[6252] <= 1'h0;
      write_done_data_log_force[6253] <= 1'h0;
      write_done_data_log_force[6254] <= 1'h0;
      write_done_data_log_force[6255] <= 1'h0;
      write_done_data_log_force[6256] <= 1'h0;
      write_done_data_log_force[6257] <= 1'h0;
      write_done_data_log_force[6258] <= 1'h0;
      write_done_data_log_force[6259] <= 1'h0;
      write_done_data_log_force[6260] <= 1'h0;
      write_done_data_log_force[6261] <= 1'h0;
      write_done_data_log_force[6262] <= 1'h0;
      write_done_data_log_force[6263] <= 1'h0;
      write_done_data_log_force[6264] <= 1'h0;
      write_done_data_log_force[6265] <= 1'h0;
      write_done_data_log_force[6266] <= 1'h0;
      write_done_data_log_force[6267] <= 1'h0;
      write_done_data_log_force[6268] <= 1'h0;
      write_done_data_log_force[6269] <= 1'h0;
      write_done_data_log_force[6270] <= 1'h0;
      write_done_data_log_force[6271] <= 1'h0;
      write_done_data_log_force[6272] <= 1'h0;
      write_done_data_log_force[6273] <= 1'h0;
      write_done_data_log_force[6274] <= 1'h0;
      write_done_data_log_force[6275] <= 1'h0;
      write_done_data_log_force[6276] <= 1'h0;
      write_done_data_log_force[6277] <= 1'h0;
      write_done_data_log_force[6278] <= 1'h0;
      write_done_data_log_force[6279] <= 1'h0;
      write_done_data_log_force[6280] <= 1'h0;
      write_done_data_log_force[6281] <= 1'h0;
      write_done_data_log_force[6282] <= 1'h0;
      write_done_data_log_force[6283] <= 1'h0;
      write_done_data_log_force[6284] <= 1'h0;
      write_done_data_log_force[6285] <= 1'h0;
      write_done_data_log_force[6286] <= 1'h0;
      write_done_data_log_force[6287] <= 1'h0;
      write_done_data_log_force[6288] <= 1'h0;
      write_done_data_log_force[6289] <= 1'h0;
      write_done_data_log_force[6290] <= 1'h0;
      write_done_data_log_force[6291] <= 1'h0;
      write_done_data_log_force[6292] <= 1'h0;
      write_done_data_log_force[6293] <= 1'h0;
      write_done_data_log_force[6294] <= 1'h0;
      write_done_data_log_force[6295] <= 1'h0;
      write_done_data_log_force[6296] <= 1'h0;
      write_done_data_log_force[6297] <= 1'h0;
      write_done_data_log_force[6298] <= 1'h0;
      write_done_data_log_force[6299] <= 1'h0;
      write_done_data_log_force[6300] <= 1'h0;
      write_done_data_log_force[6301] <= 1'h0;
      write_done_data_log_force[6302] <= 1'h0;
      write_done_data_log_force[6303] <= 1'h0;
      write_done_data_log_force[6304] <= 1'h0;
      write_done_data_log_force[6305] <= 1'h0;
      write_done_data_log_force[6306] <= 1'h0;
      write_done_data_log_force[6307] <= 1'h0;
      write_done_data_log_force[6308] <= 1'h0;
      write_done_data_log_force[6309] <= 1'h0;
      write_done_data_log_force[6310] <= 1'h0;
      write_done_data_log_force[6311] <= 1'h0;
      write_done_data_log_force[6312] <= 1'h0;
      write_done_data_log_force[6313] <= 1'h0;
      write_done_data_log_force[6314] <= 1'h0;
      write_done_data_log_force[6315] <= 1'h0;
      write_done_data_log_force[6316] <= 1'h0;
      write_done_data_log_force[6317] <= 1'h0;
      write_done_data_log_force[6318] <= 1'h0;
      write_done_data_log_force[6319] <= 1'h0;
      write_done_data_log_force[6320] <= 1'h0;
      write_done_data_log_force[6321] <= 1'h0;
      write_done_data_log_force[6322] <= 1'h0;
      write_done_data_log_force[6323] <= 1'h0;
      write_done_data_log_force[6324] <= 1'h0;
      write_done_data_log_force[6325] <= 1'h0;
      write_done_data_log_force[6326] <= 1'h0;
      write_done_data_log_force[6327] <= 1'h0;
      write_done_data_log_force[6328] <= 1'h0;
      write_done_data_log_force[6329] <= 1'h0;
      write_done_data_log_force[6330] <= 1'h0;
      write_done_data_log_force[6331] <= 1'h0;
      write_done_data_log_force[6332] <= 1'h0;
      write_done_data_log_force[6333] <= 1'h0;
      write_done_data_log_force[6334] <= 1'h0;
      write_done_data_log_force[6335] <= 1'h0;
      write_done_data_log_force[6336] <= 1'h0;
      write_done_data_log_force[6337] <= 1'h0;
      write_done_data_log_force[6338] <= 1'h0;
      write_done_data_log_force[6339] <= 1'h0;
      write_done_data_log_force[6340] <= 1'h0;
      write_done_data_log_force[6341] <= 1'h0;
      write_done_data_log_force[6342] <= 1'h0;
      write_done_data_log_force[6343] <= 1'h0;
      write_done_data_log_force[6344] <= 1'h0;
      write_done_data_log_force[6345] <= 1'h0;
      write_done_data_log_force[6346] <= 1'h0;
      write_done_data_log_force[6347] <= 1'h0;
      write_done_data_log_force[6348] <= 1'h0;
      write_done_data_log_force[6349] <= 1'h0;
      write_done_data_log_force[6350] <= 1'h0;
      write_done_data_log_force[6351] <= 1'h0;
      write_done_data_log_force[6352] <= 1'h0;
      write_done_data_log_force[6353] <= 1'h0;
      write_done_data_log_force[6354] <= 1'h0;
      write_done_data_log_force[6355] <= 1'h0;
      write_done_data_log_force[6356] <= 1'h0;
      write_done_data_log_force[6357] <= 1'h0;
      write_done_data_log_force[6358] <= 1'h0;
      write_done_data_log_force[6359] <= 1'h0;
      write_done_data_log_force[6360] <= 1'h0;
      write_done_data_log_force[6361] <= 1'h0;
      write_done_data_log_force[6362] <= 1'h0;
      write_done_data_log_force[6363] <= 1'h0;
      write_done_data_log_force[6364] <= 1'h0;
      write_done_data_log_force[6365] <= 1'h0;
      write_done_data_log_force[6366] <= 1'h0;
      write_done_data_log_force[6367] <= 1'h0;
      write_done_data_log_force[6368] <= 1'h0;
      write_done_data_log_force[6369] <= 1'h0;
      write_done_data_log_force[6370] <= 1'h0;
      write_done_data_log_force[6371] <= 1'h0;
      write_done_data_log_force[6372] <= 1'h0;
      write_done_data_log_force[6373] <= 1'h0;
      write_done_data_log_force[6374] <= 1'h0;
      write_done_data_log_force[6375] <= 1'h0;
      write_done_data_log_force[6376] <= 1'h0;
      write_done_data_log_force[6377] <= 1'h0;
      write_done_data_log_force[6378] <= 1'h0;
      write_done_data_log_force[6379] <= 1'h0;
      write_done_data_log_force[6380] <= 1'h0;
      write_done_data_log_force[6381] <= 1'h0;
      write_done_data_log_force[6382] <= 1'h0;
      write_done_data_log_force[6383] <= 1'h0;
      write_done_data_log_force[6384] <= 1'h0;
      write_done_data_log_force[6385] <= 1'h0;
      write_done_data_log_force[6386] <= 1'h0;
      write_done_data_log_force[6387] <= 1'h0;
      write_done_data_log_force[6388] <= 1'h0;
      write_done_data_log_force[6389] <= 1'h0;
      write_done_data_log_force[6390] <= 1'h0;
      write_done_data_log_force[6391] <= 1'h0;
      write_done_data_log_force[6392] <= 1'h0;
      write_done_data_log_force[6393] <= 1'h0;
      write_done_data_log_force[6394] <= 1'h0;
      write_done_data_log_force[6395] <= 1'h0;
      write_done_data_log_force[6396] <= 1'h0;
      write_done_data_log_force[6397] <= 1'h0;
      write_done_data_log_force[6398] <= 1'h0;
      write_done_data_log_force[6399] <= 1'h0;
      write_done_data_log_force[6400] <= 1'h0;
      write_done_data_log_force[6401] <= 1'h0;
      write_done_data_log_force[6402] <= 1'h0;
      write_done_data_log_force[6403] <= 1'h0;
      write_done_data_log_force[6404] <= 1'h0;
      write_done_data_log_force[6405] <= 1'h0;
      write_done_data_log_force[6406] <= 1'h0;
      write_done_data_log_force[6407] <= 1'h0;
      write_done_data_log_force[6408] <= 1'h0;
      write_done_data_log_force[6409] <= 1'h0;
      write_done_data_log_force[6410] <= 1'h0;
      write_done_data_log_force[6411] <= 1'h0;
      write_done_data_log_force[6412] <= 1'h0;
      write_done_data_log_force[6413] <= 1'h0;
      write_done_data_log_force[6414] <= 1'h0;
      write_done_data_log_force[6415] <= 1'h0;
      write_done_data_log_force[6416] <= 1'h0;
      write_done_data_log_force[6417] <= 1'h0;
      write_done_data_log_force[6418] <= 1'h0;
      write_done_data_log_force[6419] <= 1'h0;
      write_done_data_log_force[6420] <= 1'h0;
      write_done_data_log_force[6421] <= 1'h0;
      write_done_data_log_force[6422] <= 1'h0;
      write_done_data_log_force[6423] <= 1'h0;
      write_done_data_log_force[6424] <= 1'h0;
      write_done_data_log_force[6425] <= 1'h0;
      write_done_data_log_force[6426] <= 1'h0;
      write_done_data_log_force[6427] <= 1'h0;
      write_done_data_log_force[6428] <= 1'h0;
      write_done_data_log_force[6429] <= 1'h0;
      write_done_data_log_force[6430] <= 1'h0;
      write_done_data_log_force[6431] <= 1'h0;
      write_done_data_log_force[6432] <= 1'h0;
      write_done_data_log_force[6433] <= 1'h0;
      write_done_data_log_force[6434] <= 1'h0;
      write_done_data_log_force[6435] <= 1'h0;
      write_done_data_log_force[6436] <= 1'h0;
      write_done_data_log_force[6437] <= 1'h0;
      write_done_data_log_force[6438] <= 1'h0;
      write_done_data_log_force[6439] <= 1'h0;
      write_done_data_log_force[6440] <= 1'h0;
      write_done_data_log_force[6441] <= 1'h0;
      write_done_data_log_force[6442] <= 1'h0;
      write_done_data_log_force[6443] <= 1'h0;
      write_done_data_log_force[6444] <= 1'h0;
      write_done_data_log_force[6445] <= 1'h0;
      write_done_data_log_force[6446] <= 1'h0;
      write_done_data_log_force[6447] <= 1'h0;
      write_done_data_log_force[6448] <= 1'h0;
      write_done_data_log_force[6449] <= 1'h0;
      write_done_data_log_force[6450] <= 1'h0;
      write_done_data_log_force[6451] <= 1'h0;
      write_done_data_log_force[6452] <= 1'h0;
      write_done_data_log_force[6453] <= 1'h0;
      write_done_data_log_force[6454] <= 1'h0;
      write_done_data_log_force[6455] <= 1'h0;
      write_done_data_log_force[6456] <= 1'h0;
      write_done_data_log_force[6457] <= 1'h0;
      write_done_data_log_force[6458] <= 1'h0;
      write_done_data_log_force[6459] <= 1'h0;
      write_done_data_log_force[6460] <= 1'h0;
      write_done_data_log_force[6461] <= 1'h0;
      write_done_data_log_force[6462] <= 1'h0;
      write_done_data_log_force[6463] <= 1'h0;
      write_done_data_log_force[6464] <= 1'h0;
      write_done_data_log_force[6465] <= 1'h0;
      write_done_data_log_force[6466] <= 1'h0;
      write_done_data_log_force[6467] <= 1'h0;
      write_done_data_log_force[6468] <= 1'h0;
      write_done_data_log_force[6469] <= 1'h0;
      write_done_data_log_force[6470] <= 1'h0;
      write_done_data_log_force[6471] <= 1'h0;
      write_done_data_log_force[6472] <= 1'h0;
      write_done_data_log_force[6473] <= 1'h0;
      write_done_data_log_force[6474] <= 1'h0;
      write_done_data_log_force[6475] <= 1'h0;
      write_done_data_log_force[6476] <= 1'h0;
      write_done_data_log_force[6477] <= 1'h0;
      write_done_data_log_force[6478] <= 1'h0;
      write_done_data_log_force[6479] <= 1'h0;
      write_done_data_log_force[6480] <= 1'h0;
      write_done_data_log_force[6481] <= 1'h0;
      write_done_data_log_force[6482] <= 1'h0;
      write_done_data_log_force[6483] <= 1'h0;
      write_done_data_log_force[6484] <= 1'h0;
      write_done_data_log_force[6485] <= 1'h0;
      write_done_data_log_force[6486] <= 1'h0;
      write_done_data_log_force[6487] <= 1'h0;
      write_done_data_log_force[6488] <= 1'h0;
      write_done_data_log_force[6489] <= 1'h0;
      write_done_data_log_force[6490] <= 1'h0;
      write_done_data_log_force[6491] <= 1'h0;
      write_done_data_log_force[6492] <= 1'h0;
      write_done_data_log_force[6493] <= 1'h0;
      write_done_data_log_force[6494] <= 1'h0;
      write_done_data_log_force[6495] <= 1'h0;
      write_done_data_log_force[6496] <= 1'h0;
      write_done_data_log_force[6497] <= 1'h0;
      write_done_data_log_force[6498] <= 1'h0;
      write_done_data_log_force[6499] <= 1'h0;
      write_done_data_log_force[6500] <= 1'h0;
      write_done_data_log_force[6501] <= 1'h0;
      write_done_data_log_force[6502] <= 1'h0;
      write_done_data_log_force[6503] <= 1'h0;
      write_done_data_log_force[6504] <= 1'h0;
      write_done_data_log_force[6505] <= 1'h0;
      write_done_data_log_force[6506] <= 1'h0;
      write_done_data_log_force[6507] <= 1'h0;
      write_done_data_log_force[6508] <= 1'h0;
      write_done_data_log_force[6509] <= 1'h0;
      write_done_data_log_force[6510] <= 1'h0;
      write_done_data_log_force[6511] <= 1'h0;
      write_done_data_log_force[6512] <= 1'h0;
      write_done_data_log_force[6513] <= 1'h0;
      write_done_data_log_force[6514] <= 1'h0;
      write_done_data_log_force[6515] <= 1'h0;
      write_done_data_log_force[6516] <= 1'h0;
      write_done_data_log_force[6517] <= 1'h0;
      write_done_data_log_force[6518] <= 1'h0;
      write_done_data_log_force[6519] <= 1'h0;
      write_done_data_log_force[6520] <= 1'h0;
      write_done_data_log_force[6521] <= 1'h0;
      write_done_data_log_force[6522] <= 1'h0;
      write_done_data_log_force[6523] <= 1'h0;
      write_done_data_log_force[6524] <= 1'h0;
      write_done_data_log_force[6525] <= 1'h0;
      write_done_data_log_force[6526] <= 1'h0;
      write_done_data_log_force[6527] <= 1'h0;
      write_done_data_log_force[6528] <= 1'h0;
      write_done_data_log_force[6529] <= 1'h0;
      write_done_data_log_force[6530] <= 1'h0;
      write_done_data_log_force[6531] <= 1'h0;
      write_done_data_log_force[6532] <= 1'h0;
      write_done_data_log_force[6533] <= 1'h0;
      write_done_data_log_force[6534] <= 1'h0;
      write_done_data_log_force[6535] <= 1'h0;
      write_done_data_log_force[6536] <= 1'h0;
      write_done_data_log_force[6537] <= 1'h0;
      write_done_data_log_force[6538] <= 1'h0;
      write_done_data_log_force[6539] <= 1'h0;
      write_done_data_log_force[6540] <= 1'h0;
      write_done_data_log_force[6541] <= 1'h0;
      write_done_data_log_force[6542] <= 1'h0;
      write_done_data_log_force[6543] <= 1'h0;
      write_done_data_log_force[6544] <= 1'h0;
      write_done_data_log_force[6545] <= 1'h0;
      write_done_data_log_force[6546] <= 1'h0;
      write_done_data_log_force[6547] <= 1'h0;
      write_done_data_log_force[6548] <= 1'h0;
      write_done_data_log_force[6549] <= 1'h0;
      write_done_data_log_force[6550] <= 1'h0;
      write_done_data_log_force[6551] <= 1'h0;
      write_done_data_log_force[6552] <= 1'h0;
      write_done_data_log_force[6553] <= 1'h0;
      write_done_data_log_force[6554] <= 1'h0;
      write_done_data_log_force[6555] <= 1'h0;
      write_done_data_log_force[6556] <= 1'h0;
      write_done_data_log_force[6557] <= 1'h0;
      write_done_data_log_force[6558] <= 1'h0;
      write_done_data_log_force[6559] <= 1'h0;
      write_done_data_log_force[6560] <= 1'h0;
      write_done_data_log_force[6561] <= 1'h0;
      write_done_data_log_force[6562] <= 1'h0;
      write_done_data_log_force[6563] <= 1'h0;
      write_done_data_log_force[6564] <= 1'h0;
      write_done_data_log_force[6565] <= 1'h0;
      write_done_data_log_force[6566] <= 1'h0;
      write_done_data_log_force[6567] <= 1'h0;
      write_done_data_log_force[6568] <= 1'h0;
      write_done_data_log_force[6569] <= 1'h0;
      write_done_data_log_force[6570] <= 1'h0;
      write_done_data_log_force[6571] <= 1'h0;
      write_done_data_log_force[6572] <= 1'h0;
      write_done_data_log_force[6573] <= 1'h0;
      write_done_data_log_force[6574] <= 1'h0;
      write_done_data_log_force[6575] <= 1'h0;
      write_done_data_log_force[6576] <= 1'h0;
      write_done_data_log_force[6577] <= 1'h0;
      write_done_data_log_force[6578] <= 1'h0;
      write_done_data_log_force[6579] <= 1'h0;
      write_done_data_log_force[6580] <= 1'h0;
      write_done_data_log_force[6581] <= 1'h0;
      write_done_data_log_force[6582] <= 1'h0;
      write_done_data_log_force[6583] <= 1'h0;
      write_done_data_log_force[6584] <= 1'h0;
      write_done_data_log_force[6585] <= 1'h0;
      write_done_data_log_force[6586] <= 1'h0;
      write_done_data_log_force[6587] <= 1'h0;
      write_done_data_log_force[6588] <= 1'h0;
      write_done_data_log_force[6589] <= 1'h0;
      write_done_data_log_force[6590] <= 1'h0;
      write_done_data_log_force[6591] <= 1'h0;
      write_done_data_log_force[6592] <= 1'h0;
      write_done_data_log_force[6593] <= 1'h0;
      write_done_data_log_force[6594] <= 1'h0;
      write_done_data_log_force[6595] <= 1'h0;
      write_done_data_log_force[6596] <= 1'h0;
      write_done_data_log_force[6597] <= 1'h0;
      write_done_data_log_force[6598] <= 1'h0;
      write_done_data_log_force[6599] <= 1'h0;
      write_done_data_log_force[6600] <= 1'h0;
      write_done_data_log_force[6601] <= 1'h0;
      write_done_data_log_force[6602] <= 1'h0;
      write_done_data_log_force[6603] <= 1'h0;
      write_done_data_log_force[6604] <= 1'h0;
      write_done_data_log_force[6605] <= 1'h0;
      write_done_data_log_force[6606] <= 1'h0;
      write_done_data_log_force[6607] <= 1'h0;
      write_done_data_log_force[6608] <= 1'h0;
      write_done_data_log_force[6609] <= 1'h0;
      write_done_data_log_force[6610] <= 1'h0;
      write_done_data_log_force[6611] <= 1'h0;
      write_done_data_log_force[6612] <= 1'h0;
      write_done_data_log_force[6613] <= 1'h0;
      write_done_data_log_force[6614] <= 1'h0;
      write_done_data_log_force[6615] <= 1'h0;
      write_done_data_log_force[6616] <= 1'h0;
      write_done_data_log_force[6617] <= 1'h0;
      write_done_data_log_force[6618] <= 1'h0;
      write_done_data_log_force[6619] <= 1'h0;
      write_done_data_log_force[6620] <= 1'h0;
      write_done_data_log_force[6621] <= 1'h0;
      write_done_data_log_force[6622] <= 1'h0;
      write_done_data_log_force[6623] <= 1'h0;
      write_done_data_log_force[6624] <= 1'h0;
      write_done_data_log_force[6625] <= 1'h0;
      write_done_data_log_force[6626] <= 1'h0;
      write_done_data_log_force[6627] <= 1'h0;
      write_done_data_log_force[6628] <= 1'h0;
      write_done_data_log_force[6629] <= 1'h0;
      write_done_data_log_force[6630] <= 1'h0;
      write_done_data_log_force[6631] <= 1'h0;
      write_done_data_log_force[6632] <= 1'h0;
      write_done_data_log_force[6633] <= 1'h0;
      write_done_data_log_force[6634] <= 1'h0;
      write_done_data_log_force[6635] <= 1'h0;
      write_done_data_log_force[6636] <= 1'h0;
      write_done_data_log_force[6637] <= 1'h0;
      write_done_data_log_force[6638] <= 1'h0;
      write_done_data_log_force[6639] <= 1'h0;
      write_done_data_log_force[6640] <= 1'h0;
      write_done_data_log_force[6641] <= 1'h0;
      write_done_data_log_force[6642] <= 1'h0;
      write_done_data_log_force[6643] <= 1'h0;
      write_done_data_log_force[6644] <= 1'h0;
      write_done_data_log_force[6645] <= 1'h0;
      write_done_data_log_force[6646] <= 1'h0;
      write_done_data_log_force[6647] <= 1'h0;
      write_done_data_log_force[6648] <= 1'h0;
      write_done_data_log_force[6649] <= 1'h0;
      write_done_data_log_force[6650] <= 1'h0;
      write_done_data_log_force[6651] <= 1'h0;
      write_done_data_log_force[6652] <= 1'h0;
      write_done_data_log_force[6653] <= 1'h0;
      write_done_data_log_force[6654] <= 1'h0;
      write_done_data_log_force[6655] <= 1'h0;
      write_done_data_log_force[6656] <= 1'h0;
      write_done_data_log_force[6657] <= 1'h0;
      write_done_data_log_force[6658] <= 1'h0;
      write_done_data_log_force[6659] <= 1'h0;
      write_done_data_log_force[6660] <= 1'h0;
      write_done_data_log_force[6661] <= 1'h0;
      write_done_data_log_force[6662] <= 1'h0;
      write_done_data_log_force[6663] <= 1'h0;
      write_done_data_log_force[6664] <= 1'h0;
      write_done_data_log_force[6665] <= 1'h0;
      write_done_data_log_force[6666] <= 1'h0;
      write_done_data_log_force[6667] <= 1'h0;
      write_done_data_log_force[6668] <= 1'h0;
      write_done_data_log_force[6669] <= 1'h0;
      write_done_data_log_force[6670] <= 1'h0;
      write_done_data_log_force[6671] <= 1'h0;
      write_done_data_log_force[6672] <= 1'h0;
      write_done_data_log_force[6673] <= 1'h0;
      write_done_data_log_force[6674] <= 1'h0;
      write_done_data_log_force[6675] <= 1'h0;
      write_done_data_log_force[6676] <= 1'h0;
      write_done_data_log_force[6677] <= 1'h0;
      write_done_data_log_force[6678] <= 1'h0;
      write_done_data_log_force[6679] <= 1'h0;
      write_done_data_log_force[6680] <= 1'h0;
      write_done_data_log_force[6681] <= 1'h0;
      write_done_data_log_force[6682] <= 1'h0;
      write_done_data_log_force[6683] <= 1'h0;
      write_done_data_log_force[6684] <= 1'h0;
      write_done_data_log_force[6685] <= 1'h0;
      write_done_data_log_force[6686] <= 1'h0;
      write_done_data_log_force[6687] <= 1'h0;
      write_done_data_log_force[6688] <= 1'h0;
      write_done_data_log_force[6689] <= 1'h0;
      write_done_data_log_force[6690] <= 1'h0;
      write_done_data_log_force[6691] <= 1'h0;
      write_done_data_log_force[6692] <= 1'h0;
      write_done_data_log_force[6693] <= 1'h0;
      write_done_data_log_force[6694] <= 1'h0;
      write_done_data_log_force[6695] <= 1'h0;
      write_done_data_log_force[6696] <= 1'h0;
      write_done_data_log_force[6697] <= 1'h0;
      write_done_data_log_force[6698] <= 1'h0;
      write_done_data_log_force[6699] <= 1'h0;
      write_done_data_log_force[6700] <= 1'h0;
      write_done_data_log_force[6701] <= 1'h0;
      write_done_data_log_force[6702] <= 1'h0;
      write_done_data_log_force[6703] <= 1'h0;
      write_done_data_log_force[6704] <= 1'h0;
      write_done_data_log_force[6705] <= 1'h0;
      write_done_data_log_force[6706] <= 1'h0;
      write_done_data_log_force[6707] <= 1'h0;
      write_done_data_log_force[6708] <= 1'h0;
      write_done_data_log_force[6709] <= 1'h0;
      write_done_data_log_force[6710] <= 1'h0;
      write_done_data_log_force[6711] <= 1'h0;
      write_done_data_log_force[6712] <= 1'h0;
      write_done_data_log_force[6713] <= 1'h0;
      write_done_data_log_force[6714] <= 1'h0;
      write_done_data_log_force[6715] <= 1'h0;
      write_done_data_log_force[6716] <= 1'h0;
      write_done_data_log_force[6717] <= 1'h0;
      write_done_data_log_force[6718] <= 1'h0;
      write_done_data_log_force[6719] <= 1'h0;
      write_done_data_log_force[6720] <= 1'h0;
      write_done_data_log_force[6721] <= 1'h0;
      write_done_data_log_force[6722] <= 1'h0;
      write_done_data_log_force[6723] <= 1'h0;
      write_done_data_log_force[6724] <= 1'h0;
      write_done_data_log_force[6725] <= 1'h0;
      write_done_data_log_force[6726] <= 1'h0;
      write_done_data_log_force[6727] <= 1'h0;
      write_done_data_log_force[6728] <= 1'h0;
      write_done_data_log_force[6729] <= 1'h0;
      write_done_data_log_force[6730] <= 1'h0;
      write_done_data_log_force[6731] <= 1'h0;
      write_done_data_log_force[6732] <= 1'h0;
      write_done_data_log_force[6733] <= 1'h0;
      write_done_data_log_force[6734] <= 1'h0;
      write_done_data_log_force[6735] <= 1'h0;
      write_done_data_log_force[6736] <= 1'h0;
      write_done_data_log_force[6737] <= 1'h0;
      write_done_data_log_force[6738] <= 1'h0;
      write_done_data_log_force[6739] <= 1'h0;
      write_done_data_log_force[6740] <= 1'h0;
      write_done_data_log_force[6741] <= 1'h0;
      write_done_data_log_force[6742] <= 1'h0;
      write_done_data_log_force[6743] <= 1'h0;
      write_done_data_log_force[6744] <= 1'h0;
      write_done_data_log_force[6745] <= 1'h0;
      write_done_data_log_force[6746] <= 1'h0;
      write_done_data_log_force[6747] <= 1'h0;
      write_done_data_log_force[6748] <= 1'h0;
      write_done_data_log_force[6749] <= 1'h0;
      write_done_data_log_force[6750] <= 1'h0;
      write_done_data_log_force[6751] <= 1'h0;
      write_done_data_log_force[6752] <= 1'h0;
      write_done_data_log_force[6753] <= 1'h0;
      write_done_data_log_force[6754] <= 1'h0;
      write_done_data_log_force[6755] <= 1'h0;
      write_done_data_log_force[6756] <= 1'h0;
      write_done_data_log_force[6757] <= 1'h0;
      write_done_data_log_force[6758] <= 1'h0;
      write_done_data_log_force[6759] <= 1'h0;
      write_done_data_log_force[6760] <= 1'h0;
      write_done_data_log_force[6761] <= 1'h0;
      write_done_data_log_force[6762] <= 1'h0;
      write_done_data_log_force[6763] <= 1'h0;
      write_done_data_log_force[6764] <= 1'h0;
      write_done_data_log_force[6765] <= 1'h0;
      write_done_data_log_force[6766] <= 1'h0;
      write_done_data_log_force[6767] <= 1'h0;
      write_done_data_log_force[6768] <= 1'h0;
      write_done_data_log_force[6769] <= 1'h0;
      write_done_data_log_force[6770] <= 1'h0;
      write_done_data_log_force[6771] <= 1'h0;
      write_done_data_log_force[6772] <= 1'h0;
      write_done_data_log_force[6773] <= 1'h0;
      write_done_data_log_force[6774] <= 1'h0;
      write_done_data_log_force[6775] <= 1'h0;
      write_done_data_log_force[6776] <= 1'h0;
      write_done_data_log_force[6777] <= 1'h0;
      write_done_data_log_force[6778] <= 1'h0;
      write_done_data_log_force[6779] <= 1'h0;
      write_done_data_log_force[6780] <= 1'h0;
      write_done_data_log_force[6781] <= 1'h0;
      write_done_data_log_force[6782] <= 1'h0;
      write_done_data_log_force[6783] <= 1'h0;
      write_done_data_log_force[6784] <= 1'h0;
      write_done_data_log_force[6785] <= 1'h0;
      write_done_data_log_force[6786] <= 1'h0;
      write_done_data_log_force[6787] <= 1'h0;
      write_done_data_log_force[6788] <= 1'h0;
      write_done_data_log_force[6789] <= 1'h0;
      write_done_data_log_force[6790] <= 1'h0;
      write_done_data_log_force[6791] <= 1'h0;
      write_done_data_log_force[6792] <= 1'h0;
      write_done_data_log_force[6793] <= 1'h0;
      write_done_data_log_force[6794] <= 1'h0;
      write_done_data_log_force[6795] <= 1'h0;
      write_done_data_log_force[6796] <= 1'h0;
      write_done_data_log_force[6797] <= 1'h0;
      write_done_data_log_force[6798] <= 1'h0;
      write_done_data_log_force[6799] <= 1'h0;
      write_done_data_log_force[6800] <= 1'h0;
      write_done_data_log_force[6801] <= 1'h0;
      write_done_data_log_force[6802] <= 1'h0;
      write_done_data_log_force[6803] <= 1'h0;
      write_done_data_log_force[6804] <= 1'h0;
      write_done_data_log_force[6805] <= 1'h0;
      write_done_data_log_force[6806] <= 1'h0;
      write_done_data_log_force[6807] <= 1'h0;
      write_done_data_log_force[6808] <= 1'h0;
      write_done_data_log_force[6809] <= 1'h0;
      write_done_data_log_force[6810] <= 1'h0;
      write_done_data_log_force[6811] <= 1'h0;
      write_done_data_log_force[6812] <= 1'h0;
      write_done_data_log_force[6813] <= 1'h0;
      write_done_data_log_force[6814] <= 1'h0;
      write_done_data_log_force[6815] <= 1'h0;
      write_done_data_log_force[6816] <= 1'h0;
      write_done_data_log_force[6817] <= 1'h0;
      write_done_data_log_force[6818] <= 1'h0;
      write_done_data_log_force[6819] <= 1'h0;
      write_done_data_log_force[6820] <= 1'h0;
      write_done_data_log_force[6821] <= 1'h0;
      write_done_data_log_force[6822] <= 1'h0;
      write_done_data_log_force[6823] <= 1'h0;
      write_done_data_log_force[6824] <= 1'h0;
      write_done_data_log_force[6825] <= 1'h0;
      write_done_data_log_force[6826] <= 1'h0;
      write_done_data_log_force[6827] <= 1'h0;
      write_done_data_log_force[6828] <= 1'h0;
      write_done_data_log_force[6829] <= 1'h0;
      write_done_data_log_force[6830] <= 1'h0;
      write_done_data_log_force[6831] <= 1'h0;
      write_done_data_log_force[6832] <= 1'h0;
      write_done_data_log_force[6833] <= 1'h0;
      write_done_data_log_force[6834] <= 1'h0;
      write_done_data_log_force[6835] <= 1'h0;
      write_done_data_log_force[6836] <= 1'h0;
      write_done_data_log_force[6837] <= 1'h0;
      write_done_data_log_force[6838] <= 1'h0;
      write_done_data_log_force[6839] <= 1'h0;
      write_done_data_log_force[6840] <= 1'h0;
      write_done_data_log_force[6841] <= 1'h0;
      write_done_data_log_force[6842] <= 1'h0;
      write_done_data_log_force[6843] <= 1'h0;
      write_done_data_log_force[6844] <= 1'h0;
      write_done_data_log_force[6845] <= 1'h0;
      write_done_data_log_force[6846] <= 1'h0;
      write_done_data_log_force[6847] <= 1'h0;
      write_done_data_log_force[6848] <= 1'h0;
      write_done_data_log_force[6849] <= 1'h0;
      write_done_data_log_force[6850] <= 1'h0;
      write_done_data_log_force[6851] <= 1'h0;
      write_done_data_log_force[6852] <= 1'h0;
      write_done_data_log_force[6853] <= 1'h0;
      write_done_data_log_force[6854] <= 1'h0;
      write_done_data_log_force[6855] <= 1'h0;
      write_done_data_log_force[6856] <= 1'h0;
      write_done_data_log_force[6857] <= 1'h0;
      write_done_data_log_force[6858] <= 1'h0;
      write_done_data_log_force[6859] <= 1'h0;
      write_done_data_log_force[6860] <= 1'h0;
      write_done_data_log_force[6861] <= 1'h0;
      write_done_data_log_force[6862] <= 1'h0;
      write_done_data_log_force[6863] <= 1'h0;
      write_done_data_log_force[6864] <= 1'h0;
      write_done_data_log_force[6865] <= 1'h0;
      write_done_data_log_force[6866] <= 1'h0;
      write_done_data_log_force[6867] <= 1'h0;
      write_done_data_log_force[6868] <= 1'h0;
      write_done_data_log_force[6869] <= 1'h0;
      write_done_data_log_force[6870] <= 1'h0;
      write_done_data_log_force[6871] <= 1'h0;
      write_done_data_log_force[6872] <= 1'h0;
      write_done_data_log_force[6873] <= 1'h0;
      write_done_data_log_force[6874] <= 1'h0;
      write_done_data_log_force[6875] <= 1'h0;
      write_done_data_log_force[6876] <= 1'h0;
      write_done_data_log_force[6877] <= 1'h0;
      write_done_data_log_force[6878] <= 1'h0;
      write_done_data_log_force[6879] <= 1'h0;
      write_done_data_log_force[6880] <= 1'h0;
      write_done_data_log_force[6881] <= 1'h0;
      write_done_data_log_force[6882] <= 1'h0;
      write_done_data_log_force[6883] <= 1'h0;
      write_done_data_log_force[6884] <= 1'h0;
      write_done_data_log_force[6885] <= 1'h0;
      write_done_data_log_force[6886] <= 1'h0;
      write_done_data_log_force[6887] <= 1'h0;
      write_done_data_log_force[6888] <= 1'h0;
      write_done_data_log_force[6889] <= 1'h0;
      write_done_data_log_force[6890] <= 1'h0;
      write_done_data_log_force[6891] <= 1'h0;
      write_done_data_log_force[6892] <= 1'h0;
      write_done_data_log_force[6893] <= 1'h0;
      write_done_data_log_force[6894] <= 1'h0;
      write_done_data_log_force[6895] <= 1'h0;
      write_done_data_log_force[6896] <= 1'h0;
      write_done_data_log_force[6897] <= 1'h0;
      write_done_data_log_force[6898] <= 1'h0;
      write_done_data_log_force[6899] <= 1'h0;
      write_done_data_log_force[6900] <= 1'h0;
      write_done_data_log_force[6901] <= 1'h0;
      write_done_data_log_force[6902] <= 1'h0;
      write_done_data_log_force[6903] <= 1'h0;
      write_done_data_log_force[6904] <= 1'h0;
      write_done_data_log_force[6905] <= 1'h0;
      write_done_data_log_force[6906] <= 1'h0;
      write_done_data_log_force[6907] <= 1'h0;
      write_done_data_log_force[6908] <= 1'h0;
      write_done_data_log_force[6909] <= 1'h0;
      write_done_data_log_force[6910] <= 1'h0;
      write_done_data_log_force[6911] <= 1'h0;
      write_done_data_log_force[6912] <= 1'h0;
      write_done_data_log_force[6913] <= 1'h0;
      write_done_data_log_force[6914] <= 1'h0;
      write_done_data_log_force[6915] <= 1'h0;
      write_done_data_log_force[6916] <= 1'h0;
      write_done_data_log_force[6917] <= 1'h0;
      write_done_data_log_force[6918] <= 1'h0;
      write_done_data_log_force[6919] <= 1'h0;
      write_done_data_log_force[6920] <= 1'h0;
      write_done_data_log_force[6921] <= 1'h0;
      write_done_data_log_force[6922] <= 1'h0;
      write_done_data_log_force[6923] <= 1'h0;
      write_done_data_log_force[6924] <= 1'h0;
      write_done_data_log_force[6925] <= 1'h0;
      write_done_data_log_force[6926] <= 1'h0;
      write_done_data_log_force[6927] <= 1'h0;
      write_done_data_log_force[6928] <= 1'h0;
      write_done_data_log_force[6929] <= 1'h0;
      write_done_data_log_force[6930] <= 1'h0;
      write_done_data_log_force[6931] <= 1'h0;
      write_done_data_log_force[6932] <= 1'h0;
      write_done_data_log_force[6933] <= 1'h0;
      write_done_data_log_force[6934] <= 1'h0;
      write_done_data_log_force[6935] <= 1'h0;
      write_done_data_log_force[6936] <= 1'h0;
      write_done_data_log_force[6937] <= 1'h0;
      write_done_data_log_force[6938] <= 1'h0;
      write_done_data_log_force[6939] <= 1'h0;
      write_done_data_log_force[6940] <= 1'h0;
      write_done_data_log_force[6941] <= 1'h0;
      write_done_data_log_force[6942] <= 1'h0;
      write_done_data_log_force[6943] <= 1'h0;
      write_done_data_log_force[6944] <= 1'h0;
      write_done_data_log_force[6945] <= 1'h0;
      write_done_data_log_force[6946] <= 1'h0;
      write_done_data_log_force[6947] <= 1'h0;
      write_done_data_log_force[6948] <= 1'h0;
      write_done_data_log_force[6949] <= 1'h0;
      write_done_data_log_force[6950] <= 1'h0;
      write_done_data_log_force[6951] <= 1'h0;
      write_done_data_log_force[6952] <= 1'h0;
      write_done_data_log_force[6953] <= 1'h0;
      write_done_data_log_force[6954] <= 1'h0;
      write_done_data_log_force[6955] <= 1'h0;
      write_done_data_log_force[6956] <= 1'h0;
      write_done_data_log_force[6957] <= 1'h0;
      write_done_data_log_force[6958] <= 1'h0;
      write_done_data_log_force[6959] <= 1'h0;
      write_done_data_log_force[6960] <= 1'h0;
      write_done_data_log_force[6961] <= 1'h0;
      write_done_data_log_force[6962] <= 1'h0;
      write_done_data_log_force[6963] <= 1'h0;
      write_done_data_log_force[6964] <= 1'h0;
      write_done_data_log_force[6965] <= 1'h0;
      write_done_data_log_force[6966] <= 1'h0;
      write_done_data_log_force[6967] <= 1'h0;
      write_done_data_log_force[6968] <= 1'h0;
      write_done_data_log_force[6969] <= 1'h0;
      write_done_data_log_force[6970] <= 1'h0;
      write_done_data_log_force[6971] <= 1'h0;
      write_done_data_log_force[6972] <= 1'h0;
      write_done_data_log_force[6973] <= 1'h0;
      write_done_data_log_force[6974] <= 1'h0;
      write_done_data_log_force[6975] <= 1'h0;
      write_done_data_log_force[6976] <= 1'h0;
      write_done_data_log_force[6977] <= 1'h0;
      write_done_data_log_force[6978] <= 1'h0;
      write_done_data_log_force[6979] <= 1'h0;
      write_done_data_log_force[6980] <= 1'h0;
      write_done_data_log_force[6981] <= 1'h0;
      write_done_data_log_force[6982] <= 1'h0;
      write_done_data_log_force[6983] <= 1'h0;
      write_done_data_log_force[6984] <= 1'h0;
      write_done_data_log_force[6985] <= 1'h0;
      write_done_data_log_force[6986] <= 1'h0;
      write_done_data_log_force[6987] <= 1'h0;
      write_done_data_log_force[6988] <= 1'h0;
      write_done_data_log_force[6989] <= 1'h0;
      write_done_data_log_force[6990] <= 1'h0;
      write_done_data_log_force[6991] <= 1'h0;
      write_done_data_log_force[6992] <= 1'h0;
      write_done_data_log_force[6993] <= 1'h0;
      write_done_data_log_force[6994] <= 1'h0;
      write_done_data_log_force[6995] <= 1'h0;
      write_done_data_log_force[6996] <= 1'h0;
      write_done_data_log_force[6997] <= 1'h0;
      write_done_data_log_force[6998] <= 1'h0;
      write_done_data_log_force[6999] <= 1'h0;
      write_done_data_log_force[7000] <= 1'h0;
      write_done_data_log_force[7001] <= 1'h0;
      write_done_data_log_force[7002] <= 1'h0;
      write_done_data_log_force[7003] <= 1'h0;
      write_done_data_log_force[7004] <= 1'h0;
      write_done_data_log_force[7005] <= 1'h0;
      write_done_data_log_force[7006] <= 1'h0;
      write_done_data_log_force[7007] <= 1'h0;
      write_done_data_log_force[7008] <= 1'h0;
      write_done_data_log_force[7009] <= 1'h0;
      write_done_data_log_force[7010] <= 1'h0;
      write_done_data_log_force[7011] <= 1'h0;
      write_done_data_log_force[7012] <= 1'h0;
      write_done_data_log_force[7013] <= 1'h0;
      write_done_data_log_force[7014] <= 1'h0;
      write_done_data_log_force[7015] <= 1'h0;
      write_done_data_log_force[7016] <= 1'h0;
      write_done_data_log_force[7017] <= 1'h0;
      write_done_data_log_force[7018] <= 1'h0;
      write_done_data_log_force[7019] <= 1'h0;
      write_done_data_log_force[7020] <= 1'h0;
      write_done_data_log_force[7021] <= 1'h0;
      write_done_data_log_force[7022] <= 1'h0;
      write_done_data_log_force[7023] <= 1'h0;
      write_done_data_log_force[7024] <= 1'h0;
      write_done_data_log_force[7025] <= 1'h0;
      write_done_data_log_force[7026] <= 1'h0;
      write_done_data_log_force[7027] <= 1'h0;
      write_done_data_log_force[7028] <= 1'h0;
      write_done_data_log_force[7029] <= 1'h0;
      write_done_data_log_force[7030] <= 1'h0;
      write_done_data_log_force[7031] <= 1'h0;
      write_done_data_log_force[7032] <= 1'h0;
      write_done_data_log_force[7033] <= 1'h0;
      write_done_data_log_force[7034] <= 1'h0;
      write_done_data_log_force[7035] <= 1'h0;
      write_done_data_log_force[7036] <= 1'h0;
      write_done_data_log_force[7037] <= 1'h0;
      write_done_data_log_force[7038] <= 1'h0;
      write_done_data_log_force[7039] <= 1'h0;
      write_done_data_log_force[7040] <= 1'h0;
      write_done_data_log_force[7041] <= 1'h0;
      write_done_data_log_force[7042] <= 1'h0;
      write_done_data_log_force[7043] <= 1'h0;
      write_done_data_log_force[7044] <= 1'h0;
      write_done_data_log_force[7045] <= 1'h0;
      write_done_data_log_force[7046] <= 1'h0;
      write_done_data_log_force[7047] <= 1'h0;
      write_done_data_log_force[7048] <= 1'h0;
      write_done_data_log_force[7049] <= 1'h0;
      write_done_data_log_force[7050] <= 1'h0;
      write_done_data_log_force[7051] <= 1'h0;
      write_done_data_log_force[7052] <= 1'h0;
      write_done_data_log_force[7053] <= 1'h0;
      write_done_data_log_force[7054] <= 1'h0;
      write_done_data_log_force[7055] <= 1'h0;
      write_done_data_log_force[7056] <= 1'h0;
      write_done_data_log_force[7057] <= 1'h0;
      write_done_data_log_force[7058] <= 1'h0;
      write_done_data_log_force[7059] <= 1'h0;
      write_done_data_log_force[7060] <= 1'h0;
      write_done_data_log_force[7061] <= 1'h0;
      write_done_data_log_force[7062] <= 1'h0;
      write_done_data_log_force[7063] <= 1'h0;
      write_done_data_log_force[7064] <= 1'h0;
      write_done_data_log_force[7065] <= 1'h0;
      write_done_data_log_force[7066] <= 1'h0;
      write_done_data_log_force[7067] <= 1'h0;
      write_done_data_log_force[7068] <= 1'h0;
      write_done_data_log_force[7069] <= 1'h0;
      write_done_data_log_force[7070] <= 1'h0;
      write_done_data_log_force[7071] <= 1'h0;
      write_done_data_log_force[7072] <= 1'h0;
      write_done_data_log_force[7073] <= 1'h0;
      write_done_data_log_force[7074] <= 1'h0;
      write_done_data_log_force[7075] <= 1'h0;
      write_done_data_log_force[7076] <= 1'h0;
      write_done_data_log_force[7077] <= 1'h0;
      write_done_data_log_force[7078] <= 1'h0;
      write_done_data_log_force[7079] <= 1'h0;
      write_done_data_log_force[7080] <= 1'h0;
      write_done_data_log_force[7081] <= 1'h0;
      write_done_data_log_force[7082] <= 1'h0;
      write_done_data_log_force[7083] <= 1'h0;
      write_done_data_log_force[7084] <= 1'h0;
      write_done_data_log_force[7085] <= 1'h0;
      write_done_data_log_force[7086] <= 1'h0;
      write_done_data_log_force[7087] <= 1'h0;
      write_done_data_log_force[7088] <= 1'h0;
      write_done_data_log_force[7089] <= 1'h0;
      write_done_data_log_force[7090] <= 1'h0;
      write_done_data_log_force[7091] <= 1'h0;
      write_done_data_log_force[7092] <= 1'h0;
      write_done_data_log_force[7093] <= 1'h0;
      write_done_data_log_force[7094] <= 1'h0;
      write_done_data_log_force[7095] <= 1'h0;
      write_done_data_log_force[7096] <= 1'h0;
      write_done_data_log_force[7097] <= 1'h0;
      write_done_data_log_force[7098] <= 1'h0;
      write_done_data_log_force[7099] <= 1'h0;
      write_done_data_log_force[7100] <= 1'h0;
      write_done_data_log_force[7101] <= 1'h0;
      write_done_data_log_force[7102] <= 1'h0;
      write_done_data_log_force[7103] <= 1'h0;
      write_done_data_log_force[7104] <= 1'h0;
      write_done_data_log_force[7105] <= 1'h0;
      write_done_data_log_force[7106] <= 1'h0;
      write_done_data_log_force[7107] <= 1'h0;
      write_done_data_log_force[7108] <= 1'h0;
      write_done_data_log_force[7109] <= 1'h0;
      write_done_data_log_force[7110] <= 1'h0;
      write_done_data_log_force[7111] <= 1'h0;
      write_done_data_log_force[7112] <= 1'h0;
      write_done_data_log_force[7113] <= 1'h0;
      write_done_data_log_force[7114] <= 1'h0;
      write_done_data_log_force[7115] <= 1'h0;
      write_done_data_log_force[7116] <= 1'h0;
      write_done_data_log_force[7117] <= 1'h0;
      write_done_data_log_force[7118] <= 1'h0;
      write_done_data_log_force[7119] <= 1'h0;
      write_done_data_log_force[7120] <= 1'h0;
      write_done_data_log_force[7121] <= 1'h0;
      write_done_data_log_force[7122] <= 1'h0;
      write_done_data_log_force[7123] <= 1'h0;
      write_done_data_log_force[7124] <= 1'h0;
      write_done_data_log_force[7125] <= 1'h0;
      write_done_data_log_force[7126] <= 1'h0;
      write_done_data_log_force[7127] <= 1'h0;
      write_done_data_log_force[7128] <= 1'h0;
      write_done_data_log_force[7129] <= 1'h0;
      write_done_data_log_force[7130] <= 1'h0;
      write_done_data_log_force[7131] <= 1'h0;
      write_done_data_log_force[7132] <= 1'h0;
      write_done_data_log_force[7133] <= 1'h0;
      write_done_data_log_force[7134] <= 1'h0;
      write_done_data_log_force[7135] <= 1'h0;
      write_done_data_log_force[7136] <= 1'h0;
      write_done_data_log_force[7137] <= 1'h0;
      write_done_data_log_force[7138] <= 1'h0;
      write_done_data_log_force[7139] <= 1'h0;
      write_done_data_log_force[7140] <= 1'h0;
      write_done_data_log_force[7141] <= 1'h0;
      write_done_data_log_force[7142] <= 1'h0;
      write_done_data_log_force[7143] <= 1'h0;
      write_done_data_log_force[7144] <= 1'h0;
      write_done_data_log_force[7145] <= 1'h0;
      write_done_data_log_force[7146] <= 1'h0;
      write_done_data_log_force[7147] <= 1'h0;
      write_done_data_log_force[7148] <= 1'h0;
      write_done_data_log_force[7149] <= 1'h0;
      write_done_data_log_force[7150] <= 1'h0;
      write_done_data_log_force[7151] <= 1'h0;
      write_done_data_log_force[7152] <= 1'h0;
      write_done_data_log_force[7153] <= 1'h0;
      write_done_data_log_force[7154] <= 1'h0;
      write_done_data_log_force[7155] <= 1'h0;
      write_done_data_log_force[7156] <= 1'h0;
      write_done_data_log_force[7157] <= 1'h0;
      write_done_data_log_force[7158] <= 1'h0;
      write_done_data_log_force[7159] <= 1'h0;
      write_done_data_log_force[7160] <= 1'h0;
      write_done_data_log_force[7161] <= 1'h0;
      write_done_data_log_force[7162] <= 1'h0;
      write_done_data_log_force[7163] <= 1'h0;
      write_done_data_log_force[7164] <= 1'h0;
      write_done_data_log_force[7165] <= 1'h0;
      write_done_data_log_force[7166] <= 1'h0;
      write_done_data_log_force[7167] <= 1'h0;
      write_done_data_log_force[7168] <= 1'h0;
      write_done_data_log_force[7169] <= 1'h0;
      write_done_data_log_force[7170] <= 1'h0;
      write_done_data_log_force[7171] <= 1'h0;
      write_done_data_log_force[7172] <= 1'h0;
      write_done_data_log_force[7173] <= 1'h0;
      write_done_data_log_force[7174] <= 1'h0;
      write_done_data_log_force[7175] <= 1'h0;
      write_done_data_log_force[7176] <= 1'h0;
      write_done_data_log_force[7177] <= 1'h0;
      write_done_data_log_force[7178] <= 1'h0;
      write_done_data_log_force[7179] <= 1'h0;
      write_done_data_log_force[7180] <= 1'h0;
      write_done_data_log_force[7181] <= 1'h0;
      write_done_data_log_force[7182] <= 1'h0;
      write_done_data_log_force[7183] <= 1'h0;
      write_done_data_log_force[7184] <= 1'h0;
      write_done_data_log_force[7185] <= 1'h0;
      write_done_data_log_force[7186] <= 1'h0;
      write_done_data_log_force[7187] <= 1'h0;
      write_done_data_log_force[7188] <= 1'h0;
      write_done_data_log_force[7189] <= 1'h0;
      write_done_data_log_force[7190] <= 1'h0;
      write_done_data_log_force[7191] <= 1'h0;
      write_done_data_log_force[7192] <= 1'h0;
      write_done_data_log_force[7193] <= 1'h0;
      write_done_data_log_force[7194] <= 1'h0;
      write_done_data_log_force[7195] <= 1'h0;
      write_done_data_log_force[7196] <= 1'h0;
      write_done_data_log_force[7197] <= 1'h0;
      write_done_data_log_force[7198] <= 1'h0;
      write_done_data_log_force[7199] <= 1'h0;
      write_done_data_log_force[7200] <= 1'h0;
      write_done_data_log_force[7201] <= 1'h0;
      write_done_data_log_force[7202] <= 1'h0;
      write_done_data_log_force[7203] <= 1'h0;
      write_done_data_log_force[7204] <= 1'h0;
      write_done_data_log_force[7205] <= 1'h0;
      write_done_data_log_force[7206] <= 1'h0;
      write_done_data_log_force[7207] <= 1'h0;
      write_done_data_log_force[7208] <= 1'h0;
      write_done_data_log_force[7209] <= 1'h0;
      write_done_data_log_force[7210] <= 1'h0;
      write_done_data_log_force[7211] <= 1'h0;
      write_done_data_log_force[7212] <= 1'h0;
      write_done_data_log_force[7213] <= 1'h0;
      write_done_data_log_force[7214] <= 1'h0;
      write_done_data_log_force[7215] <= 1'h0;
      write_done_data_log_force[7216] <= 1'h0;
      write_done_data_log_force[7217] <= 1'h0;
      write_done_data_log_force[7218] <= 1'h0;
      write_done_data_log_force[7219] <= 1'h0;
      write_done_data_log_force[7220] <= 1'h0;
      write_done_data_log_force[7221] <= 1'h0;
      write_done_data_log_force[7222] <= 1'h0;
      write_done_data_log_force[7223] <= 1'h0;
      write_done_data_log_force[7224] <= 1'h0;
      write_done_data_log_force[7225] <= 1'h0;
      write_done_data_log_force[7226] <= 1'h0;
      write_done_data_log_force[7227] <= 1'h0;
      write_done_data_log_force[7228] <= 1'h0;
      write_done_data_log_force[7229] <= 1'h0;
      write_done_data_log_force[7230] <= 1'h0;
      write_done_data_log_force[7231] <= 1'h0;
      write_done_data_log_force[7232] <= 1'h0;
      write_done_data_log_force[7233] <= 1'h0;
      write_done_data_log_force[7234] <= 1'h0;
      write_done_data_log_force[7235] <= 1'h0;
      write_done_data_log_force[7236] <= 1'h0;
      write_done_data_log_force[7237] <= 1'h0;
      write_done_data_log_force[7238] <= 1'h0;
      write_done_data_log_force[7239] <= 1'h0;
      write_done_data_log_force[7240] <= 1'h0;
      write_done_data_log_force[7241] <= 1'h0;
      write_done_data_log_force[7242] <= 1'h0;
      write_done_data_log_force[7243] <= 1'h0;
      write_done_data_log_force[7244] <= 1'h0;
      write_done_data_log_force[7245] <= 1'h0;
      write_done_data_log_force[7246] <= 1'h0;
      write_done_data_log_force[7247] <= 1'h0;
      write_done_data_log_force[7248] <= 1'h0;
      write_done_data_log_force[7249] <= 1'h0;
      write_done_data_log_force[7250] <= 1'h0;
      write_done_data_log_force[7251] <= 1'h0;
      write_done_data_log_force[7252] <= 1'h0;
      write_done_data_log_force[7253] <= 1'h0;
      write_done_data_log_force[7254] <= 1'h0;
      write_done_data_log_force[7255] <= 1'h0;
      write_done_data_log_force[7256] <= 1'h0;
      write_done_data_log_force[7257] <= 1'h0;
      write_done_data_log_force[7258] <= 1'h0;
      write_done_data_log_force[7259] <= 1'h0;
      write_done_data_log_force[7260] <= 1'h0;
      write_done_data_log_force[7261] <= 1'h0;
      write_done_data_log_force[7262] <= 1'h0;
      write_done_data_log_force[7263] <= 1'h0;
      write_done_data_log_force[7264] <= 1'h0;
      write_done_data_log_force[7265] <= 1'h0;
      write_done_data_log_force[7266] <= 1'h0;
      write_done_data_log_force[7267] <= 1'h0;
      write_done_data_log_force[7268] <= 1'h0;
      write_done_data_log_force[7269] <= 1'h0;
      write_done_data_log_force[7270] <= 1'h0;
      write_done_data_log_force[7271] <= 1'h0;
      write_done_data_log_force[7272] <= 1'h0;
      write_done_data_log_force[7273] <= 1'h0;
      write_done_data_log_force[7274] <= 1'h0;
      write_done_data_log_force[7275] <= 1'h0;
      write_done_data_log_force[7276] <= 1'h0;
      write_done_data_log_force[7277] <= 1'h0;
      write_done_data_log_force[7278] <= 1'h0;
      write_done_data_log_force[7279] <= 1'h0;
      write_done_data_log_force[7280] <= 1'h0;
      write_done_data_log_force[7281] <= 1'h0;
      write_done_data_log_force[7282] <= 1'h0;
      write_done_data_log_force[7283] <= 1'h0;
      write_done_data_log_force[7284] <= 1'h0;
      write_done_data_log_force[7285] <= 1'h0;
      write_done_data_log_force[7286] <= 1'h0;
      write_done_data_log_force[7287] <= 1'h0;
      write_done_data_log_force[7288] <= 1'h0;
      write_done_data_log_force[7289] <= 1'h0;
      write_done_data_log_force[7290] <= 1'h0;
      write_done_data_log_force[7291] <= 1'h0;
      write_done_data_log_force[7292] <= 1'h0;
      write_done_data_log_force[7293] <= 1'h0;
      write_done_data_log_force[7294] <= 1'h0;
      write_done_data_log_force[7295] <= 1'h0;
      write_done_data_log_force[7296] <= 1'h0;
      write_done_data_log_force[7297] <= 1'h0;
      write_done_data_log_force[7298] <= 1'h0;
      write_done_data_log_force[7299] <= 1'h0;
      write_done_data_log_force[7300] <= 1'h0;
      write_done_data_log_force[7301] <= 1'h0;
      write_done_data_log_force[7302] <= 1'h0;
      write_done_data_log_force[7303] <= 1'h0;
      write_done_data_log_force[7304] <= 1'h0;
      write_done_data_log_force[7305] <= 1'h0;
      write_done_data_log_force[7306] <= 1'h0;
      write_done_data_log_force[7307] <= 1'h0;
      write_done_data_log_force[7308] <= 1'h0;
      write_done_data_log_force[7309] <= 1'h0;
      write_done_data_log_force[7310] <= 1'h0;
      write_done_data_log_force[7311] <= 1'h0;
      write_done_data_log_force[7312] <= 1'h0;
      write_done_data_log_force[7313] <= 1'h0;
      write_done_data_log_force[7314] <= 1'h0;
      write_done_data_log_force[7315] <= 1'h0;
      write_done_data_log_force[7316] <= 1'h0;
      write_done_data_log_force[7317] <= 1'h0;
      write_done_data_log_force[7318] <= 1'h0;
      write_done_data_log_force[7319] <= 1'h0;
      write_done_data_log_force[7320] <= 1'h0;
      write_done_data_log_force[7321] <= 1'h0;
      write_done_data_log_force[7322] <= 1'h0;
      write_done_data_log_force[7323] <= 1'h0;
      write_done_data_log_force[7324] <= 1'h0;
      write_done_data_log_force[7325] <= 1'h0;
      write_done_data_log_force[7326] <= 1'h0;
      write_done_data_log_force[7327] <= 1'h0;
      write_done_data_log_force[7328] <= 1'h0;
      write_done_data_log_force[7329] <= 1'h0;
      write_done_data_log_force[7330] <= 1'h0;
      write_done_data_log_force[7331] <= 1'h0;
      write_done_data_log_force[7332] <= 1'h0;
      write_done_data_log_force[7333] <= 1'h0;
      write_done_data_log_force[7334] <= 1'h0;
      write_done_data_log_force[7335] <= 1'h0;
      write_done_data_log_force[7336] <= 1'h0;
      write_done_data_log_force[7337] <= 1'h0;
      write_done_data_log_force[7338] <= 1'h0;
      write_done_data_log_force[7339] <= 1'h0;
      write_done_data_log_force[7340] <= 1'h0;
      write_done_data_log_force[7341] <= 1'h0;
      write_done_data_log_force[7342] <= 1'h0;
      write_done_data_log_force[7343] <= 1'h0;
      write_done_data_log_force[7344] <= 1'h0;
      write_done_data_log_force[7345] <= 1'h0;
      write_done_data_log_force[7346] <= 1'h0;
      write_done_data_log_force[7347] <= 1'h0;
      write_done_data_log_force[7348] <= 1'h0;
      write_done_data_log_force[7349] <= 1'h0;
      write_done_data_log_force[7350] <= 1'h0;
      write_done_data_log_force[7351] <= 1'h0;
      write_done_data_log_force[7352] <= 1'h0;
      write_done_data_log_force[7353] <= 1'h0;
      write_done_data_log_force[7354] <= 1'h0;
      write_done_data_log_force[7355] <= 1'h0;
      write_done_data_log_force[7356] <= 1'h0;
      write_done_data_log_force[7357] <= 1'h0;
      write_done_data_log_force[7358] <= 1'h0;
      write_done_data_log_force[7359] <= 1'h0;
      write_done_data_log_force[7360] <= 1'h0;
      write_done_data_log_force[7361] <= 1'h0;
      write_done_data_log_force[7362] <= 1'h0;
      write_done_data_log_force[7363] <= 1'h0;
      write_done_data_log_force[7364] <= 1'h0;
      write_done_data_log_force[7365] <= 1'h0;
      write_done_data_log_force[7366] <= 1'h0;
      write_done_data_log_force[7367] <= 1'h0;
      write_done_data_log_force[7368] <= 1'h0;
      write_done_data_log_force[7369] <= 1'h0;
      write_done_data_log_force[7370] <= 1'h0;
      write_done_data_log_force[7371] <= 1'h0;
      write_done_data_log_force[7372] <= 1'h0;
      write_done_data_log_force[7373] <= 1'h0;
      write_done_data_log_force[7374] <= 1'h0;
      write_done_data_log_force[7375] <= 1'h0;
      write_done_data_log_force[7376] <= 1'h0;
      write_done_data_log_force[7377] <= 1'h0;
      write_done_data_log_force[7378] <= 1'h0;
      write_done_data_log_force[7379] <= 1'h0;
      write_done_data_log_force[7380] <= 1'h0;
      write_done_data_log_force[7381] <= 1'h0;
      write_done_data_log_force[7382] <= 1'h0;
      write_done_data_log_force[7383] <= 1'h0;
      write_done_data_log_force[7384] <= 1'h0;
      write_done_data_log_force[7385] <= 1'h0;
      write_done_data_log_force[7386] <= 1'h0;
      write_done_data_log_force[7387] <= 1'h0;
      write_done_data_log_force[7388] <= 1'h0;
      write_done_data_log_force[7389] <= 1'h0;
      write_done_data_log_force[7390] <= 1'h0;
      write_done_data_log_force[7391] <= 1'h0;
      write_done_data_log_force[7392] <= 1'h0;
      write_done_data_log_force[7393] <= 1'h0;
      write_done_data_log_force[7394] <= 1'h0;
      write_done_data_log_force[7395] <= 1'h0;
      write_done_data_log_force[7396] <= 1'h0;
      write_done_data_log_force[7397] <= 1'h0;
      write_done_data_log_force[7398] <= 1'h0;
      write_done_data_log_force[7399] <= 1'h0;
      write_done_data_log_force[7400] <= 1'h0;
      write_done_data_log_force[7401] <= 1'h0;
      write_done_data_log_force[7402] <= 1'h0;
      write_done_data_log_force[7403] <= 1'h0;
      write_done_data_log_force[7404] <= 1'h0;
      write_done_data_log_force[7405] <= 1'h0;
      write_done_data_log_force[7406] <= 1'h0;
      write_done_data_log_force[7407] <= 1'h0;
      write_done_data_log_force[7408] <= 1'h0;
      write_done_data_log_force[7409] <= 1'h0;
      write_done_data_log_force[7410] <= 1'h0;
      write_done_data_log_force[7411] <= 1'h0;
      write_done_data_log_force[7412] <= 1'h0;
      write_done_data_log_force[7413] <= 1'h0;
      write_done_data_log_force[7414] <= 1'h0;
      write_done_data_log_force[7415] <= 1'h0;
      write_done_data_log_force[7416] <= 1'h0;
      write_done_data_log_force[7417] <= 1'h0;
      write_done_data_log_force[7418] <= 1'h0;
      write_done_data_log_force[7419] <= 1'h0;
      write_done_data_log_force[7420] <= 1'h0;
      write_done_data_log_force[7421] <= 1'h0;
      write_done_data_log_force[7422] <= 1'h0;
      write_done_data_log_force[7423] <= 1'h0;
      write_done_data_log_force[7424] <= 1'h0;
      write_done_data_log_force[7425] <= 1'h0;
      write_done_data_log_force[7426] <= 1'h0;
      write_done_data_log_force[7427] <= 1'h0;
      write_done_data_log_force[7428] <= 1'h0;
      write_done_data_log_force[7429] <= 1'h0;
      write_done_data_log_force[7430] <= 1'h0;
      write_done_data_log_force[7431] <= 1'h0;
      write_done_data_log_force[7432] <= 1'h0;
      write_done_data_log_force[7433] <= 1'h0;
      write_done_data_log_force[7434] <= 1'h0;
      write_done_data_log_force[7435] <= 1'h0;
      write_done_data_log_force[7436] <= 1'h0;
      write_done_data_log_force[7437] <= 1'h0;
      write_done_data_log_force[7438] <= 1'h0;
      write_done_data_log_force[7439] <= 1'h0;
      write_done_data_log_force[7440] <= 1'h0;
      write_done_data_log_force[7441] <= 1'h0;
      write_done_data_log_force[7442] <= 1'h0;
      write_done_data_log_force[7443] <= 1'h0;
      write_done_data_log_force[7444] <= 1'h0;
      write_done_data_log_force[7445] <= 1'h0;
      write_done_data_log_force[7446] <= 1'h0;
      write_done_data_log_force[7447] <= 1'h0;
      write_done_data_log_force[7448] <= 1'h0;
      write_done_data_log_force[7449] <= 1'h0;
      write_done_data_log_force[7450] <= 1'h0;
      write_done_data_log_force[7451] <= 1'h0;
      write_done_data_log_force[7452] <= 1'h0;
      write_done_data_log_force[7453] <= 1'h0;
      write_done_data_log_force[7454] <= 1'h0;
      write_done_data_log_force[7455] <= 1'h0;
      write_done_data_log_force[7456] <= 1'h0;
      write_done_data_log_force[7457] <= 1'h0;
      write_done_data_log_force[7458] <= 1'h0;
      write_done_data_log_force[7459] <= 1'h0;
      write_done_data_log_force[7460] <= 1'h0;
      write_done_data_log_force[7461] <= 1'h0;
      write_done_data_log_force[7462] <= 1'h0;
      write_done_data_log_force[7463] <= 1'h0;
      write_done_data_log_force[7464] <= 1'h0;
      write_done_data_log_force[7465] <= 1'h0;
      write_done_data_log_force[7466] <= 1'h0;
      write_done_data_log_force[7467] <= 1'h0;
      write_done_data_log_force[7468] <= 1'h0;
      write_done_data_log_force[7469] <= 1'h0;
      write_done_data_log_force[7470] <= 1'h0;
      write_done_data_log_force[7471] <= 1'h0;
      write_done_data_log_force[7472] <= 1'h0;
      write_done_data_log_force[7473] <= 1'h0;
      write_done_data_log_force[7474] <= 1'h0;
      write_done_data_log_force[7475] <= 1'h0;
      write_done_data_log_force[7476] <= 1'h0;
      write_done_data_log_force[7477] <= 1'h0;
      write_done_data_log_force[7478] <= 1'h0;
      write_done_data_log_force[7479] <= 1'h0;
      write_done_data_log_force[7480] <= 1'h0;
      write_done_data_log_force[7481] <= 1'h0;
      write_done_data_log_force[7482] <= 1'h0;
      write_done_data_log_force[7483] <= 1'h0;
      write_done_data_log_force[7484] <= 1'h0;
      write_done_data_log_force[7485] <= 1'h0;
      write_done_data_log_force[7486] <= 1'h0;
      write_done_data_log_force[7487] <= 1'h0;
      write_done_data_log_force[7488] <= 1'h0;
      write_done_data_log_force[7489] <= 1'h0;
      write_done_data_log_force[7490] <= 1'h0;
      write_done_data_log_force[7491] <= 1'h0;
      write_done_data_log_force[7492] <= 1'h0;
      write_done_data_log_force[7493] <= 1'h0;
      write_done_data_log_force[7494] <= 1'h0;
      write_done_data_log_force[7495] <= 1'h0;
      write_done_data_log_force[7496] <= 1'h0;
      write_done_data_log_force[7497] <= 1'h0;
      write_done_data_log_force[7498] <= 1'h0;
      write_done_data_log_force[7499] <= 1'h0;
      write_done_data_log_force[7500] <= 1'h0;
      write_done_data_log_force[7501] <= 1'h0;
      write_done_data_log_force[7502] <= 1'h0;
      write_done_data_log_force[7503] <= 1'h0;
      write_done_data_log_force[7504] <= 1'h0;
      write_done_data_log_force[7505] <= 1'h0;
      write_done_data_log_force[7506] <= 1'h0;
      write_done_data_log_force[7507] <= 1'h0;
      write_done_data_log_force[7508] <= 1'h0;
      write_done_data_log_force[7509] <= 1'h0;
      write_done_data_log_force[7510] <= 1'h0;
      write_done_data_log_force[7511] <= 1'h0;
      write_done_data_log_force[7512] <= 1'h0;
      write_done_data_log_force[7513] <= 1'h0;
      write_done_data_log_force[7514] <= 1'h0;
      write_done_data_log_force[7515] <= 1'h0;
      write_done_data_log_force[7516] <= 1'h0;
      write_done_data_log_force[7517] <= 1'h0;
      write_done_data_log_force[7518] <= 1'h0;
      write_done_data_log_force[7519] <= 1'h0;
      write_done_data_log_force[7520] <= 1'h0;
      write_done_data_log_force[7521] <= 1'h0;
      write_done_data_log_force[7522] <= 1'h0;
      write_done_data_log_force[7523] <= 1'h0;
      write_done_data_log_force[7524] <= 1'h0;
      write_done_data_log_force[7525] <= 1'h0;
      write_done_data_log_force[7526] <= 1'h0;
      write_done_data_log_force[7527] <= 1'h0;
      write_done_data_log_force[7528] <= 1'h0;
      write_done_data_log_force[7529] <= 1'h0;
      write_done_data_log_force[7530] <= 1'h0;
      write_done_data_log_force[7531] <= 1'h0;
      write_done_data_log_force[7532] <= 1'h0;
      write_done_data_log_force[7533] <= 1'h0;
      write_done_data_log_force[7534] <= 1'h0;
      write_done_data_log_force[7535] <= 1'h0;
      write_done_data_log_force[7536] <= 1'h0;
      write_done_data_log_force[7537] <= 1'h0;
      write_done_data_log_force[7538] <= 1'h0;
      write_done_data_log_force[7539] <= 1'h0;
      write_done_data_log_force[7540] <= 1'h0;
      write_done_data_log_force[7541] <= 1'h0;
      write_done_data_log_force[7542] <= 1'h0;
      write_done_data_log_force[7543] <= 1'h0;
      write_done_data_log_force[7544] <= 1'h0;
      write_done_data_log_force[7545] <= 1'h0;
      write_done_data_log_force[7546] <= 1'h0;
      write_done_data_log_force[7547] <= 1'h0;
      write_done_data_log_force[7548] <= 1'h0;
      write_done_data_log_force[7549] <= 1'h0;
      write_done_data_log_force[7550] <= 1'h0;
      write_done_data_log_force[7551] <= 1'h0;
      write_done_data_log_force[7552] <= 1'h0;
      write_done_data_log_force[7553] <= 1'h0;
      write_done_data_log_force[7554] <= 1'h0;
      write_done_data_log_force[7555] <= 1'h0;
      write_done_data_log_force[7556] <= 1'h0;
      write_done_data_log_force[7557] <= 1'h0;
      write_done_data_log_force[7558] <= 1'h0;
      write_done_data_log_force[7559] <= 1'h0;
      write_done_data_log_force[7560] <= 1'h0;
      write_done_data_log_force[7561] <= 1'h0;
      write_done_data_log_force[7562] <= 1'h0;
      write_done_data_log_force[7563] <= 1'h0;
      write_done_data_log_force[7564] <= 1'h0;
      write_done_data_log_force[7565] <= 1'h0;
      write_done_data_log_force[7566] <= 1'h0;
      write_done_data_log_force[7567] <= 1'h0;
      write_done_data_log_force[7568] <= 1'h0;
      write_done_data_log_force[7569] <= 1'h0;
      write_done_data_log_force[7570] <= 1'h0;
      write_done_data_log_force[7571] <= 1'h0;
      write_done_data_log_force[7572] <= 1'h0;
      write_done_data_log_force[7573] <= 1'h0;
      write_done_data_log_force[7574] <= 1'h0;
      write_done_data_log_force[7575] <= 1'h0;
      write_done_data_log_force[7576] <= 1'h0;
      write_done_data_log_force[7577] <= 1'h0;
      write_done_data_log_force[7578] <= 1'h0;
      write_done_data_log_force[7579] <= 1'h0;
      write_done_data_log_force[7580] <= 1'h0;
      write_done_data_log_force[7581] <= 1'h0;
      write_done_data_log_force[7582] <= 1'h0;
      write_done_data_log_force[7583] <= 1'h0;
      write_done_data_log_force[7584] <= 1'h0;
      write_done_data_log_force[7585] <= 1'h0;
      write_done_data_log_force[7586] <= 1'h0;
      write_done_data_log_force[7587] <= 1'h0;
      write_done_data_log_force[7588] <= 1'h0;
      write_done_data_log_force[7589] <= 1'h0;
      write_done_data_log_force[7590] <= 1'h0;
      write_done_data_log_force[7591] <= 1'h0;
      write_done_data_log_force[7592] <= 1'h0;
      write_done_data_log_force[7593] <= 1'h0;
      write_done_data_log_force[7594] <= 1'h0;
      write_done_data_log_force[7595] <= 1'h0;
      write_done_data_log_force[7596] <= 1'h0;
      write_done_data_log_force[7597] <= 1'h0;
      write_done_data_log_force[7598] <= 1'h0;
      write_done_data_log_force[7599] <= 1'h0;
      write_done_data_log_force[7600] <= 1'h0;
      write_done_data_log_force[7601] <= 1'h0;
      write_done_data_log_force[7602] <= 1'h0;
      write_done_data_log_force[7603] <= 1'h0;
      write_done_data_log_force[7604] <= 1'h0;
      write_done_data_log_force[7605] <= 1'h0;
      write_done_data_log_force[7606] <= 1'h0;
      write_done_data_log_force[7607] <= 1'h0;
      write_done_data_log_force[7608] <= 1'h0;
      write_done_data_log_force[7609] <= 1'h0;
      write_done_data_log_force[7610] <= 1'h0;
      write_done_data_log_force[7611] <= 1'h0;
      write_done_data_log_force[7612] <= 1'h0;
      write_done_data_log_force[7613] <= 1'h0;
      write_done_data_log_force[7614] <= 1'h0;
      write_done_data_log_force[7615] <= 1'h0;
      write_done_data_log_force[7616] <= 1'h0;
      write_done_data_log_force[7617] <= 1'h0;
      write_done_data_log_force[7618] <= 1'h0;
      write_done_data_log_force[7619] <= 1'h0;
      write_done_data_log_force[7620] <= 1'h0;
      write_done_data_log_force[7621] <= 1'h0;
      write_done_data_log_force[7622] <= 1'h0;
      write_done_data_log_force[7623] <= 1'h0;
      write_done_data_log_force[7624] <= 1'h0;
      write_done_data_log_force[7625] <= 1'h0;
      write_done_data_log_force[7626] <= 1'h0;
      write_done_data_log_force[7627] <= 1'h0;
      write_done_data_log_force[7628] <= 1'h0;
      write_done_data_log_force[7629] <= 1'h0;
      write_done_data_log_force[7630] <= 1'h0;
      write_done_data_log_force[7631] <= 1'h0;
      write_done_data_log_force[7632] <= 1'h0;
      write_done_data_log_force[7633] <= 1'h0;
      write_done_data_log_force[7634] <= 1'h0;
      write_done_data_log_force[7635] <= 1'h0;
      write_done_data_log_force[7636] <= 1'h0;
      write_done_data_log_force[7637] <= 1'h0;
      write_done_data_log_force[7638] <= 1'h0;
      write_done_data_log_force[7639] <= 1'h0;
      write_done_data_log_force[7640] <= 1'h0;
      write_done_data_log_force[7641] <= 1'h0;
      write_done_data_log_force[7642] <= 1'h0;
      write_done_data_log_force[7643] <= 1'h0;
      write_done_data_log_force[7644] <= 1'h0;
      write_done_data_log_force[7645] <= 1'h0;
      write_done_data_log_force[7646] <= 1'h0;
      write_done_data_log_force[7647] <= 1'h0;
      write_done_data_log_force[7648] <= 1'h0;
      write_done_data_log_force[7649] <= 1'h0;
      write_done_data_log_force[7650] <= 1'h0;
      write_done_data_log_force[7651] <= 1'h0;
      write_done_data_log_force[7652] <= 1'h0;
      write_done_data_log_force[7653] <= 1'h0;
      write_done_data_log_force[7654] <= 1'h0;
      write_done_data_log_force[7655] <= 1'h0;
      write_done_data_log_force[7656] <= 1'h0;
      write_done_data_log_force[7657] <= 1'h0;
      write_done_data_log_force[7658] <= 1'h0;
      write_done_data_log_force[7659] <= 1'h0;
      write_done_data_log_force[7660] <= 1'h0;
      write_done_data_log_force[7661] <= 1'h0;
      write_done_data_log_force[7662] <= 1'h0;
      write_done_data_log_force[7663] <= 1'h0;
      write_done_data_log_force[7664] <= 1'h0;
      write_done_data_log_force[7665] <= 1'h0;
      write_done_data_log_force[7666] <= 1'h0;
      write_done_data_log_force[7667] <= 1'h0;
      write_done_data_log_force[7668] <= 1'h0;
      write_done_data_log_force[7669] <= 1'h0;
      write_done_data_log_force[7670] <= 1'h0;
      write_done_data_log_force[7671] <= 1'h0;
      write_done_data_log_force[7672] <= 1'h0;
      write_done_data_log_force[7673] <= 1'h0;
      write_done_data_log_force[7674] <= 1'h0;
      write_done_data_log_force[7675] <= 1'h0;
      write_done_data_log_force[7676] <= 1'h0;
      write_done_data_log_force[7677] <= 1'h0;
      write_done_data_log_force[7678] <= 1'h0;
      write_done_data_log_force[7679] <= 1'h0;
      write_done_data_log_force[7680] <= 1'h0;
      write_done_data_log_force[7681] <= 1'h0;
      write_done_data_log_force[7682] <= 1'h0;
      write_done_data_log_force[7683] <= 1'h0;
      write_done_data_log_force[7684] <= 1'h0;
      write_done_data_log_force[7685] <= 1'h0;
      write_done_data_log_force[7686] <= 1'h0;
      write_done_data_log_force[7687] <= 1'h0;
      write_done_data_log_force[7688] <= 1'h0;
      write_done_data_log_force[7689] <= 1'h0;
      write_done_data_log_force[7690] <= 1'h0;
      write_done_data_log_force[7691] <= 1'h0;
      write_done_data_log_force[7692] <= 1'h0;
      write_done_data_log_force[7693] <= 1'h0;
      write_done_data_log_force[7694] <= 1'h0;
      write_done_data_log_force[7695] <= 1'h0;
      write_done_data_log_force[7696] <= 1'h0;
      write_done_data_log_force[7697] <= 1'h0;
      write_done_data_log_force[7698] <= 1'h0;
      write_done_data_log_force[7699] <= 1'h0;
      write_done_data_log_force[7700] <= 1'h0;
      write_done_data_log_force[7701] <= 1'h0;
      write_done_data_log_force[7702] <= 1'h0;
      write_done_data_log_force[7703] <= 1'h0;
      write_done_data_log_force[7704] <= 1'h0;
      write_done_data_log_force[7705] <= 1'h0;
      write_done_data_log_force[7706] <= 1'h0;
      write_done_data_log_force[7707] <= 1'h0;
      write_done_data_log_force[7708] <= 1'h0;
      write_done_data_log_force[7709] <= 1'h0;
      write_done_data_log_force[7710] <= 1'h0;
      write_done_data_log_force[7711] <= 1'h0;
      write_done_data_log_force[7712] <= 1'h0;
      write_done_data_log_force[7713] <= 1'h0;
      write_done_data_log_force[7714] <= 1'h0;
      write_done_data_log_force[7715] <= 1'h0;
      write_done_data_log_force[7716] <= 1'h0;
      write_done_data_log_force[7717] <= 1'h0;
      write_done_data_log_force[7718] <= 1'h0;
      write_done_data_log_force[7719] <= 1'h0;
      write_done_data_log_force[7720] <= 1'h0;
      write_done_data_log_force[7721] <= 1'h0;
      write_done_data_log_force[7722] <= 1'h0;
      write_done_data_log_force[7723] <= 1'h0;
      write_done_data_log_force[7724] <= 1'h0;
      write_done_data_log_force[7725] <= 1'h0;
      write_done_data_log_force[7726] <= 1'h0;
      write_done_data_log_force[7727] <= 1'h0;
      write_done_data_log_force[7728] <= 1'h0;
      write_done_data_log_force[7729] <= 1'h0;
      write_done_data_log_force[7730] <= 1'h0;
      write_done_data_log_force[7731] <= 1'h0;
      write_done_data_log_force[7732] <= 1'h0;
      write_done_data_log_force[7733] <= 1'h0;
      write_done_data_log_force[7734] <= 1'h0;
      write_done_data_log_force[7735] <= 1'h0;
      write_done_data_log_force[7736] <= 1'h0;
      write_done_data_log_force[7737] <= 1'h0;
      write_done_data_log_force[7738] <= 1'h0;
      write_done_data_log_force[7739] <= 1'h0;
      write_done_data_log_force[7740] <= 1'h0;
      write_done_data_log_force[7741] <= 1'h0;
      write_done_data_log_force[7742] <= 1'h0;
      write_done_data_log_force[7743] <= 1'h0;
      write_done_data_log_force[7744] <= 1'h0;
      write_done_data_log_force[7745] <= 1'h0;
      write_done_data_log_force[7746] <= 1'h0;
      write_done_data_log_force[7747] <= 1'h0;
      write_done_data_log_force[7748] <= 1'h0;
      write_done_data_log_force[7749] <= 1'h0;
      write_done_data_log_force[7750] <= 1'h0;
      write_done_data_log_force[7751] <= 1'h0;
      write_done_data_log_force[7752] <= 1'h0;
      write_done_data_log_force[7753] <= 1'h0;
      write_done_data_log_force[7754] <= 1'h0;
      write_done_data_log_force[7755] <= 1'h0;
      write_done_data_log_force[7756] <= 1'h0;
      write_done_data_log_force[7757] <= 1'h0;
      write_done_data_log_force[7758] <= 1'h0;
      write_done_data_log_force[7759] <= 1'h0;
      write_done_data_log_force[7760] <= 1'h0;
      write_done_data_log_force[7761] <= 1'h0;
      write_done_data_log_force[7762] <= 1'h0;
      write_done_data_log_force[7763] <= 1'h0;
      write_done_data_log_force[7764] <= 1'h0;
      write_done_data_log_force[7765] <= 1'h0;
      write_done_data_log_force[7766] <= 1'h0;
      write_done_data_log_force[7767] <= 1'h0;
      write_done_data_log_force[7768] <= 1'h0;
      write_done_data_log_force[7769] <= 1'h0;
      write_done_data_log_force[7770] <= 1'h0;
      write_done_data_log_force[7771] <= 1'h0;
      write_done_data_log_force[7772] <= 1'h0;
      write_done_data_log_force[7773] <= 1'h0;
      write_done_data_log_force[7774] <= 1'h0;
      write_done_data_log_force[7775] <= 1'h0;
      write_done_data_log_force[7776] <= 1'h0;
      write_done_data_log_force[7777] <= 1'h0;
      write_done_data_log_force[7778] <= 1'h0;
      write_done_data_log_force[7779] <= 1'h0;
      write_done_data_log_force[7780] <= 1'h0;
      write_done_data_log_force[7781] <= 1'h0;
      write_done_data_log_force[7782] <= 1'h0;
      write_done_data_log_force[7783] <= 1'h0;
      write_done_data_log_force[7784] <= 1'h0;
      write_done_data_log_force[7785] <= 1'h0;
      write_done_data_log_force[7786] <= 1'h0;
      write_done_data_log_force[7787] <= 1'h0;
      write_done_data_log_force[7788] <= 1'h0;
      write_done_data_log_force[7789] <= 1'h0;
      write_done_data_log_force[7790] <= 1'h0;
      write_done_data_log_force[7791] <= 1'h0;
      write_done_data_log_force[7792] <= 1'h0;
      write_done_data_log_force[7793] <= 1'h0;
      write_done_data_log_force[7794] <= 1'h0;
      write_done_data_log_force[7795] <= 1'h0;
      write_done_data_log_force[7796] <= 1'h0;
      write_done_data_log_force[7797] <= 1'h0;
      write_done_data_log_force[7798] <= 1'h0;
      write_done_data_log_force[7799] <= 1'h0;
      write_done_data_log_force[7800] <= 1'h0;
      write_done_data_log_force[7801] <= 1'h0;
      write_done_data_log_force[7802] <= 1'h0;
      write_done_data_log_force[7803] <= 1'h0;
      write_done_data_log_force[7804] <= 1'h0;
      write_done_data_log_force[7805] <= 1'h0;
      write_done_data_log_force[7806] <= 1'h0;
      write_done_data_log_force[7807] <= 1'h0;
      write_done_data_log_force[7808] <= 1'h0;
      write_done_data_log_force[7809] <= 1'h0;
      write_done_data_log_force[7810] <= 1'h0;
      write_done_data_log_force[7811] <= 1'h0;
      write_done_data_log_force[7812] <= 1'h0;
      write_done_data_log_force[7813] <= 1'h0;
      write_done_data_log_force[7814] <= 1'h0;
      write_done_data_log_force[7815] <= 1'h0;
      write_done_data_log_force[7816] <= 1'h0;
      write_done_data_log_force[7817] <= 1'h0;
      write_done_data_log_force[7818] <= 1'h0;
      write_done_data_log_force[7819] <= 1'h0;
      write_done_data_log_force[7820] <= 1'h0;
      write_done_data_log_force[7821] <= 1'h0;
      write_done_data_log_force[7822] <= 1'h0;
      write_done_data_log_force[7823] <= 1'h0;
      write_done_data_log_force[7824] <= 1'h0;
      write_done_data_log_force[7825] <= 1'h0;
      write_done_data_log_force[7826] <= 1'h0;
      write_done_data_log_force[7827] <= 1'h0;
      write_done_data_log_force[7828] <= 1'h0;
      write_done_data_log_force[7829] <= 1'h0;
      write_done_data_log_force[7830] <= 1'h0;
      write_done_data_log_force[7831] <= 1'h0;
      write_done_data_log_force[7832] <= 1'h0;
      write_done_data_log_force[7833] <= 1'h0;
      write_done_data_log_force[7834] <= 1'h0;
      write_done_data_log_force[7835] <= 1'h0;
      write_done_data_log_force[7836] <= 1'h0;
      write_done_data_log_force[7837] <= 1'h0;
      write_done_data_log_force[7838] <= 1'h0;
      write_done_data_log_force[7839] <= 1'h0;
      write_done_data_log_force[7840] <= 1'h0;
      write_done_data_log_force[7841] <= 1'h0;
      write_done_data_log_force[7842] <= 1'h0;
      write_done_data_log_force[7843] <= 1'h0;
      write_done_data_log_force[7844] <= 1'h0;
      write_done_data_log_force[7845] <= 1'h0;
      write_done_data_log_force[7846] <= 1'h0;
      write_done_data_log_force[7847] <= 1'h0;
      write_done_data_log_force[7848] <= 1'h0;
      write_done_data_log_force[7849] <= 1'h0;
      write_done_data_log_force[7850] <= 1'h0;
      write_done_data_log_force[7851] <= 1'h0;
      write_done_data_log_force[7852] <= 1'h0;
      write_done_data_log_force[7853] <= 1'h0;
      write_done_data_log_force[7854] <= 1'h0;
      write_done_data_log_force[7855] <= 1'h0;
      write_done_data_log_force[7856] <= 1'h0;
      write_done_data_log_force[7857] <= 1'h0;
      write_done_data_log_force[7858] <= 1'h0;
      write_done_data_log_force[7859] <= 1'h0;
      write_done_data_log_force[7860] <= 1'h0;
      write_done_data_log_force[7861] <= 1'h0;
      write_done_data_log_force[7862] <= 1'h0;
      write_done_data_log_force[7863] <= 1'h0;
      write_done_data_log_force[7864] <= 1'h0;
      write_done_data_log_force[7865] <= 1'h0;
      write_done_data_log_force[7866] <= 1'h0;
      write_done_data_log_force[7867] <= 1'h0;
      write_done_data_log_force[7868] <= 1'h0;
      write_done_data_log_force[7869] <= 1'h0;
      write_done_data_log_force[7870] <= 1'h0;
      write_done_data_log_force[7871] <= 1'h0;
      write_done_data_log_force[7872] <= 1'h0;
      write_done_data_log_force[7873] <= 1'h0;
      write_done_data_log_force[7874] <= 1'h0;
      write_done_data_log_force[7875] <= 1'h0;
      write_done_data_log_force[7876] <= 1'h0;
      write_done_data_log_force[7877] <= 1'h0;
      write_done_data_log_force[7878] <= 1'h0;
      write_done_data_log_force[7879] <= 1'h0;
      write_done_data_log_force[7880] <= 1'h0;
      write_done_data_log_force[7881] <= 1'h0;
      write_done_data_log_force[7882] <= 1'h0;
      write_done_data_log_force[7883] <= 1'h0;
      write_done_data_log_force[7884] <= 1'h0;
      write_done_data_log_force[7885] <= 1'h0;
      write_done_data_log_force[7886] <= 1'h0;
      write_done_data_log_force[7887] <= 1'h0;
      write_done_data_log_force[7888] <= 1'h0;
      write_done_data_log_force[7889] <= 1'h0;
      write_done_data_log_force[7890] <= 1'h0;
      write_done_data_log_force[7891] <= 1'h0;
      write_done_data_log_force[7892] <= 1'h0;
      write_done_data_log_force[7893] <= 1'h0;
      write_done_data_log_force[7894] <= 1'h0;
      write_done_data_log_force[7895] <= 1'h0;
      write_done_data_log_force[7896] <= 1'h0;
      write_done_data_log_force[7897] <= 1'h0;
      write_done_data_log_force[7898] <= 1'h0;
      write_done_data_log_force[7899] <= 1'h0;
      write_done_data_log_force[7900] <= 1'h0;
      write_done_data_log_force[7901] <= 1'h0;
      write_done_data_log_force[7902] <= 1'h0;
      write_done_data_log_force[7903] <= 1'h0;
      write_done_data_log_force[7904] <= 1'h0;
      write_done_data_log_force[7905] <= 1'h0;
      write_done_data_log_force[7906] <= 1'h0;
      write_done_data_log_force[7907] <= 1'h0;
      write_done_data_log_force[7908] <= 1'h0;
      write_done_data_log_force[7909] <= 1'h0;
      write_done_data_log_force[7910] <= 1'h0;
      write_done_data_log_force[7911] <= 1'h0;
      write_done_data_log_force[7912] <= 1'h0;
      write_done_data_log_force[7913] <= 1'h0;
      write_done_data_log_force[7914] <= 1'h0;
      write_done_data_log_force[7915] <= 1'h0;
      write_done_data_log_force[7916] <= 1'h0;
      write_done_data_log_force[7917] <= 1'h0;
      write_done_data_log_force[7918] <= 1'h0;
      write_done_data_log_force[7919] <= 1'h0;
      write_done_data_log_force[7920] <= 1'h0;
      write_done_data_log_force[7921] <= 1'h0;
      write_done_data_log_force[7922] <= 1'h0;
      write_done_data_log_force[7923] <= 1'h0;
      write_done_data_log_force[7924] <= 1'h0;
      write_done_data_log_force[7925] <= 1'h0;
      write_done_data_log_force[7926] <= 1'h0;
      write_done_data_log_force[7927] <= 1'h0;
      write_done_data_log_force[7928] <= 1'h0;
      write_done_data_log_force[7929] <= 1'h0;
      write_done_data_log_force[7930] <= 1'h0;
      write_done_data_log_force[7931] <= 1'h0;
      write_done_data_log_force[7932] <= 1'h0;
      write_done_data_log_force[7933] <= 1'h0;
      write_done_data_log_force[7934] <= 1'h0;
      write_done_data_log_force[7935] <= 1'h0;
      write_done_data_log_force[7936] <= 1'h0;
      write_done_data_log_force[7937] <= 1'h0;
      write_done_data_log_force[7938] <= 1'h0;
      write_done_data_log_force[7939] <= 1'h0;
      write_done_data_log_force[7940] <= 1'h0;
      write_done_data_log_force[7941] <= 1'h0;
      write_done_data_log_force[7942] <= 1'h0;
      write_done_data_log_force[7943] <= 1'h0;
      write_done_data_log_force[7944] <= 1'h0;
      write_done_data_log_force[7945] <= 1'h0;
      write_done_data_log_force[7946] <= 1'h0;
      write_done_data_log_force[7947] <= 1'h0;
      write_done_data_log_force[7948] <= 1'h0;
      write_done_data_log_force[7949] <= 1'h0;
      write_done_data_log_force[7950] <= 1'h0;
      write_done_data_log_force[7951] <= 1'h0;
      write_done_data_log_force[7952] <= 1'h0;
      write_done_data_log_force[7953] <= 1'h0;
      write_done_data_log_force[7954] <= 1'h0;
      write_done_data_log_force[7955] <= 1'h0;
      write_done_data_log_force[7956] <= 1'h0;
      write_done_data_log_force[7957] <= 1'h0;
      write_done_data_log_force[7958] <= 1'h0;
      write_done_data_log_force[7959] <= 1'h0;
      write_done_data_log_force[7960] <= 1'h0;
      write_done_data_log_force[7961] <= 1'h0;
      write_done_data_log_force[7962] <= 1'h0;
      write_done_data_log_force[7963] <= 1'h0;
      write_done_data_log_force[7964] <= 1'h0;
      write_done_data_log_force[7965] <= 1'h0;
      write_done_data_log_force[7966] <= 1'h0;
      write_done_data_log_force[7967] <= 1'h0;
      write_done_data_log_force[7968] <= 1'h0;
      write_done_data_log_force[7969] <= 1'h0;
      write_done_data_log_force[7970] <= 1'h0;
      write_done_data_log_force[7971] <= 1'h0;
      write_done_data_log_force[7972] <= 1'h0;
      write_done_data_log_force[7973] <= 1'h0;
      write_done_data_log_force[7974] <= 1'h0;
      write_done_data_log_force[7975] <= 1'h0;
      write_done_data_log_force[7976] <= 1'h0;
      write_done_data_log_force[7977] <= 1'h0;
      write_done_data_log_force[7978] <= 1'h0;
      write_done_data_log_force[7979] <= 1'h0;
      write_done_data_log_force[7980] <= 1'h0;
      write_done_data_log_force[7981] <= 1'h0;
      write_done_data_log_force[7982] <= 1'h0;
      write_done_data_log_force[7983] <= 1'h0;
      write_done_data_log_force[7984] <= 1'h0;
      write_done_data_log_force[7985] <= 1'h0;
      write_done_data_log_force[7986] <= 1'h0;
      write_done_data_log_force[7987] <= 1'h0;
      write_done_data_log_force[7988] <= 1'h0;
      write_done_data_log_force[7989] <= 1'h0;
      write_done_data_log_force[7990] <= 1'h0;
      write_done_data_log_force[7991] <= 1'h0;
      write_done_data_log_force[7992] <= 1'h0;
      write_done_data_log_force[7993] <= 1'h0;
      write_done_data_log_force[7994] <= 1'h0;
      write_done_data_log_force[7995] <= 1'h0;
      write_done_data_log_force[7996] <= 1'h0;
      write_done_data_log_force[7997] <= 1'h0;
      write_done_data_log_force[7998] <= 1'h0;
      write_done_data_log_force[7999] <= 1'h0;
      write_done_data_log_force[8000] <= 1'h0;
      write_done_data_log_force[8001] <= 1'h0;
      write_done_data_log_force[8002] <= 1'h0;
      write_done_data_log_force[8003] <= 1'h0;
      write_done_data_log_force[8004] <= 1'h0;
      write_done_data_log_force[8005] <= 1'h0;
      write_done_data_log_force[8006] <= 1'h0;
      write_done_data_log_force[8007] <= 1'h0;
      write_done_data_log_force[8008] <= 1'h0;
      write_done_data_log_force[8009] <= 1'h0;
      write_done_data_log_force[8010] <= 1'h0;
      write_done_data_log_force[8011] <= 1'h0;
      write_done_data_log_force[8012] <= 1'h0;
      write_done_data_log_force[8013] <= 1'h0;
      write_done_data_log_force[8014] <= 1'h0;
      write_done_data_log_force[8015] <= 1'h0;
      write_done_data_log_force[8016] <= 1'h0;
      write_done_data_log_force[8017] <= 1'h0;
      write_done_data_log_force[8018] <= 1'h0;
      write_done_data_log_force[8019] <= 1'h0;
      write_done_data_log_force[8020] <= 1'h0;
      write_done_data_log_force[8021] <= 1'h0;
      write_done_data_log_force[8022] <= 1'h0;
      write_done_data_log_force[8023] <= 1'h0;
      write_done_data_log_force[8024] <= 1'h0;
      write_done_data_log_force[8025] <= 1'h0;
      write_done_data_log_force[8026] <= 1'h0;
      write_done_data_log_force[8027] <= 1'h0;
      write_done_data_log_force[8028] <= 1'h0;
      write_done_data_log_force[8029] <= 1'h0;
      write_done_data_log_force[8030] <= 1'h0;
      write_done_data_log_force[8031] <= 1'h0;
      write_done_data_log_force[8032] <= 1'h0;
      write_done_data_log_force[8033] <= 1'h0;
      write_done_data_log_force[8034] <= 1'h0;
      write_done_data_log_force[8035] <= 1'h0;
      write_done_data_log_force[8036] <= 1'h0;
      write_done_data_log_force[8037] <= 1'h0;
      write_done_data_log_force[8038] <= 1'h0;
      write_done_data_log_force[8039] <= 1'h0;
      write_done_data_log_force[8040] <= 1'h0;
      write_done_data_log_force[8041] <= 1'h0;
      write_done_data_log_force[8042] <= 1'h0;
      write_done_data_log_force[8043] <= 1'h0;
      write_done_data_log_force[8044] <= 1'h0;
      write_done_data_log_force[8045] <= 1'h0;
      write_done_data_log_force[8046] <= 1'h0;
      write_done_data_log_force[8047] <= 1'h0;
      write_done_data_log_force[8048] <= 1'h0;
      write_done_data_log_force[8049] <= 1'h0;
      write_done_data_log_force[8050] <= 1'h0;
      write_done_data_log_force[8051] <= 1'h0;
      write_done_data_log_force[8052] <= 1'h0;
      write_done_data_log_force[8053] <= 1'h0;
      write_done_data_log_force[8054] <= 1'h0;
      write_done_data_log_force[8055] <= 1'h0;
      write_done_data_log_force[8056] <= 1'h0;
      write_done_data_log_force[8057] <= 1'h0;
      write_done_data_log_force[8058] <= 1'h0;
      write_done_data_log_force[8059] <= 1'h0;
      write_done_data_log_force[8060] <= 1'h0;
      write_done_data_log_force[8061] <= 1'h0;
      write_done_data_log_force[8062] <= 1'h0;
      write_done_data_log_force[8063] <= 1'h0;
      write_done_data_log_force[8064] <= 1'h0;
      write_done_data_log_force[8065] <= 1'h0;
      write_done_data_log_force[8066] <= 1'h0;
      write_done_data_log_force[8067] <= 1'h0;
      write_done_data_log_force[8068] <= 1'h0;
      write_done_data_log_force[8069] <= 1'h0;
      write_done_data_log_force[8070] <= 1'h0;
      write_done_data_log_force[8071] <= 1'h0;
      write_done_data_log_force[8072] <= 1'h0;
      write_done_data_log_force[8073] <= 1'h0;
      write_done_data_log_force[8074] <= 1'h0;
      write_done_data_log_force[8075] <= 1'h0;
      write_done_data_log_force[8076] <= 1'h0;
      write_done_data_log_force[8077] <= 1'h0;
      write_done_data_log_force[8078] <= 1'h0;
      write_done_data_log_force[8079] <= 1'h0;
      write_done_data_log_force[8080] <= 1'h0;
      write_done_data_log_force[8081] <= 1'h0;
      write_done_data_log_force[8082] <= 1'h0;
      write_done_data_log_force[8083] <= 1'h0;
      write_done_data_log_force[8084] <= 1'h0;
      write_done_data_log_force[8085] <= 1'h0;
      write_done_data_log_force[8086] <= 1'h0;
      write_done_data_log_force[8087] <= 1'h0;
      write_done_data_log_force[8088] <= 1'h0;
      write_done_data_log_force[8089] <= 1'h0;
      write_done_data_log_force[8090] <= 1'h0;
      write_done_data_log_force[8091] <= 1'h0;
      write_done_data_log_force[8092] <= 1'h0;
      write_done_data_log_force[8093] <= 1'h0;
      write_done_data_log_force[8094] <= 1'h0;
      write_done_data_log_force[8095] <= 1'h0;
      write_done_data_log_force[8096] <= 1'h0;
      write_done_data_log_force[8097] <= 1'h0;
      write_done_data_log_force[8098] <= 1'h0;
      write_done_data_log_force[8099] <= 1'h0;
      write_done_data_log_force[8100] <= 1'h0;
      write_done_data_log_force[8101] <= 1'h0;
      write_done_data_log_force[8102] <= 1'h0;
      write_done_data_log_force[8103] <= 1'h0;
      write_done_data_log_force[8104] <= 1'h0;
      write_done_data_log_force[8105] <= 1'h0;
      write_done_data_log_force[8106] <= 1'h0;
      write_done_data_log_force[8107] <= 1'h0;
      write_done_data_log_force[8108] <= 1'h0;
      write_done_data_log_force[8109] <= 1'h0;
      write_done_data_log_force[8110] <= 1'h0;
      write_done_data_log_force[8111] <= 1'h0;
      write_done_data_log_force[8112] <= 1'h0;
      write_done_data_log_force[8113] <= 1'h0;
      write_done_data_log_force[8114] <= 1'h0;
      write_done_data_log_force[8115] <= 1'h0;
      write_done_data_log_force[8116] <= 1'h0;
      write_done_data_log_force[8117] <= 1'h0;
      write_done_data_log_force[8118] <= 1'h0;
      write_done_data_log_force[8119] <= 1'h0;
      write_done_data_log_force[8120] <= 1'h0;
      write_done_data_log_force[8121] <= 1'h0;
      write_done_data_log_force[8122] <= 1'h0;
      write_done_data_log_force[8123] <= 1'h0;
      write_done_data_log_force[8124] <= 1'h0;
      write_done_data_log_force[8125] <= 1'h0;
      write_done_data_log_force[8126] <= 1'h0;
      write_done_data_log_force[8127] <= 1'h0;
      write_done_data_log_force[8128] <= 1'h0;
      write_done_data_log_force[8129] <= 1'h0;
      write_done_data_log_force[8130] <= 1'h0;
      write_done_data_log_force[8131] <= 1'h0;
      write_done_data_log_force[8132] <= 1'h0;
      write_done_data_log_force[8133] <= 1'h0;
      write_done_data_log_force[8134] <= 1'h0;
      write_done_data_log_force[8135] <= 1'h0;
      write_done_data_log_force[8136] <= 1'h0;
      write_done_data_log_force[8137] <= 1'h0;
      write_done_data_log_force[8138] <= 1'h0;
      write_done_data_log_force[8139] <= 1'h0;
      write_done_data_log_force[8140] <= 1'h0;
      write_done_data_log_force[8141] <= 1'h0;
      write_done_data_log_force[8142] <= 1'h0;
      write_done_data_log_force[8143] <= 1'h0;
      write_done_data_log_force[8144] <= 1'h0;
      write_done_data_log_force[8145] <= 1'h0;
      write_done_data_log_force[8146] <= 1'h0;
      write_done_data_log_force[8147] <= 1'h0;
      write_done_data_log_force[8148] <= 1'h0;
      write_done_data_log_force[8149] <= 1'h0;
      write_done_data_log_force[8150] <= 1'h0;
      write_done_data_log_force[8151] <= 1'h0;
      write_done_data_log_force[8152] <= 1'h0;
      write_done_data_log_force[8153] <= 1'h0;
      write_done_data_log_force[8154] <= 1'h0;
      write_done_data_log_force[8155] <= 1'h0;
      write_done_data_log_force[8156] <= 1'h0;
      write_done_data_log_force[8157] <= 1'h0;
      write_done_data_log_force[8158] <= 1'h0;
      write_done_data_log_force[8159] <= 1'h0;
      write_done_data_log_force[8160] <= 1'h0;
      write_done_data_log_force[8161] <= 1'h0;
      write_done_data_log_force[8162] <= 1'h0;
      write_done_data_log_force[8163] <= 1'h0;
      write_done_data_log_force[8164] <= 1'h0;
      write_done_data_log_force[8165] <= 1'h0;
      write_done_data_log_force[8166] <= 1'h0;
      write_done_data_log_force[8167] <= 1'h0;
      write_done_data_log_force[8168] <= 1'h0;
      write_done_data_log_force[8169] <= 1'h0;
      write_done_data_log_force[8170] <= 1'h0;
      write_done_data_log_force[8171] <= 1'h0;
      write_done_data_log_force[8172] <= 1'h0;
      write_done_data_log_force[8173] <= 1'h0;
      write_done_data_log_force[8174] <= 1'h0;
      write_done_data_log_force[8175] <= 1'h0;
      write_done_data_log_force[8176] <= 1'h0;
      write_done_data_log_force[8177] <= 1'h0;
      write_done_data_log_force[8178] <= 1'h0;
      write_done_data_log_force[8179] <= 1'h0;
      write_done_data_log_force[8180] <= 1'h0;
      write_done_data_log_force[8181] <= 1'h0;
      write_done_data_log_force[8182] <= 1'h0;
      write_done_data_log_force[8183] <= 1'h0;
      write_done_data_log_force[8184] <= 1'h0;
      write_done_data_log_force[8185] <= 1'h0;
      write_done_data_log_force[8186] <= 1'h0;
      write_done_data_log_force[8187] <= 1'h0;
      write_done_data_log_force[8188] <= 1'h0;
      write_done_data_log_force[8189] <= 1'h0;
      write_done_data_log_force[8190] <= 1'h0;
      write_done_data_log_force[8191] <= 1'h0;
      write_done_data_log_force[8192] <= 1'h0;
      write_done_data_log_force[8193] <= 1'h0;
      write_done_data_log_force[8194] <= 1'h0;
      write_done_data_log_force[8195] <= 1'h0;
      write_done_data_log_force[8196] <= 1'h0;
      write_done_data_log_force[8197] <= 1'h0;
      write_done_data_log_force[8198] <= 1'h0;
      write_done_data_log_force[8199] <= 1'h0;
      write_done_data_log_force[8200] <= 1'h0;
      write_done_data_log_force[8201] <= 1'h0;
      write_done_data_log_force[8202] <= 1'h0;
      write_done_data_log_force[8203] <= 1'h0;
      write_done_data_log_force[8204] <= 1'h0;
      write_done_data_log_force[8205] <= 1'h0;
      write_done_data_log_force[8206] <= 1'h0;
      write_done_data_log_force[8207] <= 1'h0;
      write_done_data_log_force[8208] <= 1'h0;
      write_done_data_log_force[8209] <= 1'h0;
      write_done_data_log_force[8210] <= 1'h0;
      write_done_data_log_force[8211] <= 1'h0;
      write_done_data_log_force[8212] <= 1'h0;
      write_done_data_log_force[8213] <= 1'h0;
      write_done_data_log_force[8214] <= 1'h0;
      write_done_data_log_force[8215] <= 1'h0;
      write_done_data_log_force[8216] <= 1'h0;
      write_done_data_log_force[8217] <= 1'h0;
      write_done_data_log_force[8218] <= 1'h0;
      write_done_data_log_force[8219] <= 1'h0;
      write_done_data_log_force[8220] <= 1'h0;
      write_done_data_log_force[8221] <= 1'h0;
      write_done_data_log_force[8222] <= 1'h0;
      write_done_data_log_force[8223] <= 1'h0;
      write_done_data_log_force[8224] <= 1'h0;
      write_done_data_log_force[8225] <= 1'h0;
      write_done_data_log_force[8226] <= 1'h0;
      write_done_data_log_force[8227] <= 1'h0;
      write_done_data_log_force[8228] <= 1'h0;
      write_done_data_log_force[8229] <= 1'h0;
      write_done_data_log_force[8230] <= 1'h0;
      write_done_data_log_force[8231] <= 1'h0;
      write_done_data_log_force[8232] <= 1'h0;
      write_done_data_log_force[8233] <= 1'h0;
      write_done_data_log_force[8234] <= 1'h0;
      write_done_data_log_force[8235] <= 1'h0;
      write_done_data_log_force[8236] <= 1'h0;
      write_done_data_log_force[8237] <= 1'h0;
      write_done_data_log_force[8238] <= 1'h0;
      write_done_data_log_force[8239] <= 1'h0;
      write_done_data_log_force[8240] <= 1'h0;
      write_done_data_log_force[8241] <= 1'h0;
      write_done_data_log_force[8242] <= 1'h0;
      write_done_data_log_force[8243] <= 1'h0;
      write_done_data_log_force[8244] <= 1'h0;
      write_done_data_log_force[8245] <= 1'h0;
      write_done_data_log_force[8246] <= 1'h0;
      write_done_data_log_force[8247] <= 1'h0;
      write_done_data_log_force[8248] <= 1'h0;
      write_done_data_log_force[8249] <= 1'h0;
      write_done_data_log_force[8250] <= 1'h0;
      write_done_data_log_force[8251] <= 1'h0;
      write_done_data_log_force[8252] <= 1'h0;
      write_done_data_log_force[8253] <= 1'h0;
      write_done_data_log_force[8254] <= 1'h0;
      write_done_data_log_force[8255] <= 1'h0;
      write_done_data_log_force[8256] <= 1'h0;
      write_done_data_log_force[8257] <= 1'h0;
      write_done_data_log_force[8258] <= 1'h0;
      write_done_data_log_force[8259] <= 1'h0;
      write_done_data_log_force[8260] <= 1'h0;
      write_done_data_log_force[8261] <= 1'h0;
      write_done_data_log_force[8262] <= 1'h0;
      write_done_data_log_force[8263] <= 1'h0;
      write_done_data_log_force[8264] <= 1'h0;
      write_done_data_log_force[8265] <= 1'h0;
      write_done_data_log_force[8266] <= 1'h0;
      write_done_data_log_force[8267] <= 1'h0;
      write_done_data_log_force[8268] <= 1'h0;
      write_done_data_log_force[8269] <= 1'h0;
      write_done_data_log_force[8270] <= 1'h0;
      write_done_data_log_force[8271] <= 1'h0;
      write_done_data_log_force[8272] <= 1'h0;
      write_done_data_log_force[8273] <= 1'h0;
      write_done_data_log_force[8274] <= 1'h0;
      write_done_data_log_force[8275] <= 1'h0;
      write_done_data_log_force[8276] <= 1'h0;
      write_done_data_log_force[8277] <= 1'h0;
      write_done_data_log_force[8278] <= 1'h0;
      write_done_data_log_force[8279] <= 1'h0;
      write_done_data_log_force[8280] <= 1'h0;
      write_done_data_log_force[8281] <= 1'h0;
      write_done_data_log_force[8282] <= 1'h0;
      write_done_data_log_force[8283] <= 1'h0;
      write_done_data_log_force[8284] <= 1'h0;
      write_done_data_log_force[8285] <= 1'h0;
      write_done_data_log_force[8286] <= 1'h0;
      write_done_data_log_force[8287] <= 1'h0;
      write_done_data_log_force[8288] <= 1'h0;
      write_done_data_log_force[8289] <= 1'h0;
      write_done_data_log_force[8290] <= 1'h0;
      write_done_data_log_force[8291] <= 1'h0;
      write_done_data_log_force[8292] <= 1'h0;
      write_done_data_log_force[8293] <= 1'h0;
      write_done_data_log_force[8294] <= 1'h0;
      write_done_data_log_force[8295] <= 1'h0;
      write_done_data_log_force[8296] <= 1'h0;
      write_done_data_log_force[8297] <= 1'h0;
      write_done_data_log_force[8298] <= 1'h0;
      write_done_data_log_force[8299] <= 1'h0;
      write_done_data_log_force[8300] <= 1'h0;
      write_done_data_log_force[8301] <= 1'h0;
      write_done_data_log_force[8302] <= 1'h0;
      write_done_data_log_force[8303] <= 1'h0;
      write_done_data_log_force[8304] <= 1'h0;
      write_done_data_log_force[8305] <= 1'h0;
      write_done_data_log_force[8306] <= 1'h0;
      write_done_data_log_force[8307] <= 1'h0;
      write_done_data_log_force[8308] <= 1'h0;
      write_done_data_log_force[8309] <= 1'h0;
      write_done_data_log_force[8310] <= 1'h0;
      write_done_data_log_force[8311] <= 1'h0;
      write_done_data_log_force[8312] <= 1'h0;
      write_done_data_log_force[8313] <= 1'h0;
      write_done_data_log_force[8314] <= 1'h0;
      write_done_data_log_force[8315] <= 1'h0;
      write_done_data_log_force[8316] <= 1'h0;
      write_done_data_log_force[8317] <= 1'h0;
      write_done_data_log_force[8318] <= 1'h0;
      write_done_data_log_force[8319] <= 1'h0;

      // Input data for write_address_data_log
      write_address_data_log_force[   0] <= 6'h00;
      write_address_data_log_force[   1] <= 6'h01;
      write_address_data_log_force[   2] <= 6'h02;
      write_address_data_log_force[   3] <= 6'h03;
      write_address_data_log_force[   4] <= 6'h04;
      write_address_data_log_force[   5] <= 6'h05;
      write_address_data_log_force[   6] <= 6'h06;
      write_address_data_log_force[   7] <= 6'h07;
      write_address_data_log_force[   8] <= 6'h08;
      write_address_data_log_force[   9] <= 6'h09;
      write_address_data_log_force[  10] <= 6'h0a;
      write_address_data_log_force[  11] <= 6'h0b;
      write_address_data_log_force[  12] <= 6'h0c;
      write_address_data_log_force[  13] <= 6'h0d;
      write_address_data_log_force[  14] <= 6'h0e;
      write_address_data_log_force[  15] <= 6'h0f;
      write_address_data_log_force[  16] <= 6'h10;
      write_address_data_log_force[  17] <= 6'h11;
      write_address_data_log_force[  18] <= 6'h12;
      write_address_data_log_force[  19] <= 6'h13;
      write_address_data_log_force[  20] <= 6'h14;
      write_address_data_log_force[  21] <= 6'h15;
      write_address_data_log_force[  22] <= 6'h16;
      write_address_data_log_force[  23] <= 6'h17;
      write_address_data_log_force[  24] <= 6'h18;
      write_address_data_log_force[  25] <= 6'h19;
      write_address_data_log_force[  26] <= 6'h1a;
      write_address_data_log_force[  27] <= 6'h1b;
      write_address_data_log_force[  28] <= 6'h1c;
      write_address_data_log_force[  29] <= 6'h1d;
      write_address_data_log_force[  30] <= 6'h1e;
      write_address_data_log_force[  31] <= 6'h1f;
      write_address_data_log_force[  32] <= 6'h20;
      write_address_data_log_force[  33] <= 6'h21;
      write_address_data_log_force[  34] <= 6'h22;
      write_address_data_log_force[  35] <= 6'h23;
      write_address_data_log_force[  36] <= 6'h24;
      write_address_data_log_force[  37] <= 6'h25;
      write_address_data_log_force[  38] <= 6'h26;
      write_address_data_log_force[  39] <= 6'h27;
      write_address_data_log_force[  40] <= 6'h28;
      write_address_data_log_force[  41] <= 6'h29;
      write_address_data_log_force[  42] <= 6'h2a;
      write_address_data_log_force[  43] <= 6'h2b;
      write_address_data_log_force[  44] <= 6'h2c;
      write_address_data_log_force[  45] <= 6'h2d;
      write_address_data_log_force[  46] <= 6'h2e;
      write_address_data_log_force[  47] <= 6'h2f;
      write_address_data_log_force[  48] <= 6'h30;
      write_address_data_log_force[  49] <= 6'h31;
      write_address_data_log_force[  50] <= 6'h32;
      write_address_data_log_force[  51] <= 6'h33;
      write_address_data_log_force[  52] <= 6'h34;
      write_address_data_log_force[  53] <= 6'h35;
      write_address_data_log_force[  54] <= 6'h36;
      write_address_data_log_force[  55] <= 6'h37;
      write_address_data_log_force[  56] <= 6'h38;
      write_address_data_log_force[  57] <= 6'h39;
      write_address_data_log_force[  58] <= 6'h3a;
      write_address_data_log_force[  59] <= 6'h3b;
      write_address_data_log_force[  60] <= 6'h3c;
      write_address_data_log_force[  61] <= 6'h3d;
      write_address_data_log_force[  62] <= 6'h3e;
      write_address_data_log_force[  63] <= 6'h3f;
      write_address_data_log_force[  64] <= 6'h00;
      write_address_data_log_force[  65] <= 6'h00;
      write_address_data_log_force[  66] <= 6'h00;
      write_address_data_log_force[  67] <= 6'h00;
      write_address_data_log_force[  68] <= 6'h00;
      write_address_data_log_force[  69] <= 6'h00;
      write_address_data_log_force[  70] <= 6'h00;
      write_address_data_log_force[  71] <= 6'h00;
      write_address_data_log_force[  72] <= 6'h00;
      write_address_data_log_force[  73] <= 6'h00;
      write_address_data_log_force[  74] <= 6'h00;
      write_address_data_log_force[  75] <= 6'h00;
      write_address_data_log_force[  76] <= 6'h00;
      write_address_data_log_force[  77] <= 6'h00;
      write_address_data_log_force[  78] <= 6'h00;
      write_address_data_log_force[  79] <= 6'h00;
      write_address_data_log_force[  80] <= 6'h00;
      write_address_data_log_force[  81] <= 6'h00;
      write_address_data_log_force[  82] <= 6'h00;
      write_address_data_log_force[  83] <= 6'h00;
      write_address_data_log_force[  84] <= 6'h00;
      write_address_data_log_force[  85] <= 6'h00;
      write_address_data_log_force[  86] <= 6'h00;
      write_address_data_log_force[  87] <= 6'h00;
      write_address_data_log_force[  88] <= 6'h00;
      write_address_data_log_force[  89] <= 6'h00;
      write_address_data_log_force[  90] <= 6'h00;
      write_address_data_log_force[  91] <= 6'h00;
      write_address_data_log_force[  92] <= 6'h00;
      write_address_data_log_force[  93] <= 6'h00;
      write_address_data_log_force[  94] <= 6'h00;
      write_address_data_log_force[  95] <= 6'h00;
      write_address_data_log_force[  96] <= 6'h00;
      write_address_data_log_force[  97] <= 6'h00;
      write_address_data_log_force[  98] <= 6'h00;
      write_address_data_log_force[  99] <= 6'h00;
      write_address_data_log_force[ 100] <= 6'h00;
      write_address_data_log_force[ 101] <= 6'h00;
      write_address_data_log_force[ 102] <= 6'h00;
      write_address_data_log_force[ 103] <= 6'h00;
      write_address_data_log_force[ 104] <= 6'h00;
      write_address_data_log_force[ 105] <= 6'h00;
      write_address_data_log_force[ 106] <= 6'h00;
      write_address_data_log_force[ 107] <= 6'h00;
      write_address_data_log_force[ 108] <= 6'h00;
      write_address_data_log_force[ 109] <= 6'h00;
      write_address_data_log_force[ 110] <= 6'h00;
      write_address_data_log_force[ 111] <= 6'h00;
      write_address_data_log_force[ 112] <= 6'h00;
      write_address_data_log_force[ 113] <= 6'h00;
      write_address_data_log_force[ 114] <= 6'h00;
      write_address_data_log_force[ 115] <= 6'h00;
      write_address_data_log_force[ 116] <= 6'h00;
      write_address_data_log_force[ 117] <= 6'h00;
      write_address_data_log_force[ 118] <= 6'h00;
      write_address_data_log_force[ 119] <= 6'h00;
      write_address_data_log_force[ 120] <= 6'h00;
      write_address_data_log_force[ 121] <= 6'h00;
      write_address_data_log_force[ 122] <= 6'h00;
      write_address_data_log_force[ 123] <= 6'h00;
      write_address_data_log_force[ 124] <= 6'h00;
      write_address_data_log_force[ 125] <= 6'h00;
      write_address_data_log_force[ 126] <= 6'h00;
      write_address_data_log_force[ 127] <= 6'h00;
      write_address_data_log_force[ 128] <= 6'h00;
      write_address_data_log_force[ 129] <= 6'h00;
      write_address_data_log_force[ 130] <= 6'h00;
      write_address_data_log_force[ 131] <= 6'h00;
      write_address_data_log_force[ 132] <= 6'h00;
      write_address_data_log_force[ 133] <= 6'h00;
      write_address_data_log_force[ 134] <= 6'h00;
      write_address_data_log_force[ 135] <= 6'h00;
      write_address_data_log_force[ 136] <= 6'h00;
      write_address_data_log_force[ 137] <= 6'h00;
      write_address_data_log_force[ 138] <= 6'h00;
      write_address_data_log_force[ 139] <= 6'h00;
      write_address_data_log_force[ 140] <= 6'h00;
      write_address_data_log_force[ 141] <= 6'h00;
      write_address_data_log_force[ 142] <= 6'h00;
      write_address_data_log_force[ 143] <= 6'h00;
      write_address_data_log_force[ 144] <= 6'h00;
      write_address_data_log_force[ 145] <= 6'h00;
      write_address_data_log_force[ 146] <= 6'h00;
      write_address_data_log_force[ 147] <= 6'h00;
      write_address_data_log_force[ 148] <= 6'h00;
      write_address_data_log_force[ 149] <= 6'h00;
      write_address_data_log_force[ 150] <= 6'h00;
      write_address_data_log_force[ 151] <= 6'h00;
      write_address_data_log_force[ 152] <= 6'h00;
      write_address_data_log_force[ 153] <= 6'h00;
      write_address_data_log_force[ 154] <= 6'h00;
      write_address_data_log_force[ 155] <= 6'h00;
      write_address_data_log_force[ 156] <= 6'h00;
      write_address_data_log_force[ 157] <= 6'h00;
      write_address_data_log_force[ 158] <= 6'h00;
      write_address_data_log_force[ 159] <= 6'h00;
      write_address_data_log_force[ 160] <= 6'h00;
      write_address_data_log_force[ 161] <= 6'h00;
      write_address_data_log_force[ 162] <= 6'h00;
      write_address_data_log_force[ 163] <= 6'h00;
      write_address_data_log_force[ 164] <= 6'h00;
      write_address_data_log_force[ 165] <= 6'h00;
      write_address_data_log_force[ 166] <= 6'h00;
      write_address_data_log_force[ 167] <= 6'h00;
      write_address_data_log_force[ 168] <= 6'h00;
      write_address_data_log_force[ 169] <= 6'h00;
      write_address_data_log_force[ 170] <= 6'h00;
      write_address_data_log_force[ 171] <= 6'h00;
      write_address_data_log_force[ 172] <= 6'h00;
      write_address_data_log_force[ 173] <= 6'h00;
      write_address_data_log_force[ 174] <= 6'h00;
      write_address_data_log_force[ 175] <= 6'h00;
      write_address_data_log_force[ 176] <= 6'h00;
      write_address_data_log_force[ 177] <= 6'h00;
      write_address_data_log_force[ 178] <= 6'h00;
      write_address_data_log_force[ 179] <= 6'h00;
      write_address_data_log_force[ 180] <= 6'h00;
      write_address_data_log_force[ 181] <= 6'h00;
      write_address_data_log_force[ 182] <= 6'h00;
      write_address_data_log_force[ 183] <= 6'h00;
      write_address_data_log_force[ 184] <= 6'h00;
      write_address_data_log_force[ 185] <= 6'h00;
      write_address_data_log_force[ 186] <= 6'h00;
      write_address_data_log_force[ 187] <= 6'h00;
      write_address_data_log_force[ 188] <= 6'h00;
      write_address_data_log_force[ 189] <= 6'h00;
      write_address_data_log_force[ 190] <= 6'h00;
      write_address_data_log_force[ 191] <= 6'h00;
      write_address_data_log_force[ 192] <= 6'h00;
      write_address_data_log_force[ 193] <= 6'h00;
      write_address_data_log_force[ 194] <= 6'h00;
      write_address_data_log_force[ 195] <= 6'h00;
      write_address_data_log_force[ 196] <= 6'h00;
      write_address_data_log_force[ 197] <= 6'h00;
      write_address_data_log_force[ 198] <= 6'h00;
      write_address_data_log_force[ 199] <= 6'h00;
      write_address_data_log_force[ 200] <= 6'h00;
      write_address_data_log_force[ 201] <= 6'h00;
      write_address_data_log_force[ 202] <= 6'h00;
      write_address_data_log_force[ 203] <= 6'h00;
      write_address_data_log_force[ 204] <= 6'h00;
      write_address_data_log_force[ 205] <= 6'h00;
      write_address_data_log_force[ 206] <= 6'h00;
      write_address_data_log_force[ 207] <= 6'h00;
      write_address_data_log_force[ 208] <= 6'h00;
      write_address_data_log_force[ 209] <= 6'h00;
      write_address_data_log_force[ 210] <= 6'h00;
      write_address_data_log_force[ 211] <= 6'h00;
      write_address_data_log_force[ 212] <= 6'h00;
      write_address_data_log_force[ 213] <= 6'h00;
      write_address_data_log_force[ 214] <= 6'h00;
      write_address_data_log_force[ 215] <= 6'h00;
      write_address_data_log_force[ 216] <= 6'h00;
      write_address_data_log_force[ 217] <= 6'h00;
      write_address_data_log_force[ 218] <= 6'h00;
      write_address_data_log_force[ 219] <= 6'h00;
      write_address_data_log_force[ 220] <= 6'h00;
      write_address_data_log_force[ 221] <= 6'h00;
      write_address_data_log_force[ 222] <= 6'h00;
      write_address_data_log_force[ 223] <= 6'h00;
      write_address_data_log_force[ 224] <= 6'h00;
      write_address_data_log_force[ 225] <= 6'h00;
      write_address_data_log_force[ 226] <= 6'h00;
      write_address_data_log_force[ 227] <= 6'h00;
      write_address_data_log_force[ 228] <= 6'h00;
      write_address_data_log_force[ 229] <= 6'h00;
      write_address_data_log_force[ 230] <= 6'h00;
      write_address_data_log_force[ 231] <= 6'h00;
      write_address_data_log_force[ 232] <= 6'h00;
      write_address_data_log_force[ 233] <= 6'h00;
      write_address_data_log_force[ 234] <= 6'h00;
      write_address_data_log_force[ 235] <= 6'h00;
      write_address_data_log_force[ 236] <= 6'h00;
      write_address_data_log_force[ 237] <= 6'h00;
      write_address_data_log_force[ 238] <= 6'h00;
      write_address_data_log_force[ 239] <= 6'h00;
      write_address_data_log_force[ 240] <= 6'h00;
      write_address_data_log_force[ 241] <= 6'h00;
      write_address_data_log_force[ 242] <= 6'h00;
      write_address_data_log_force[ 243] <= 6'h00;
      write_address_data_log_force[ 244] <= 6'h00;
      write_address_data_log_force[ 245] <= 6'h00;
      write_address_data_log_force[ 246] <= 6'h00;
      write_address_data_log_force[ 247] <= 6'h00;
      write_address_data_log_force[ 248] <= 6'h00;
      write_address_data_log_force[ 249] <= 6'h00;
      write_address_data_log_force[ 250] <= 6'h00;
      write_address_data_log_force[ 251] <= 6'h00;
      write_address_data_log_force[ 252] <= 6'h00;
      write_address_data_log_force[ 253] <= 6'h00;
      write_address_data_log_force[ 254] <= 6'h00;
      write_address_data_log_force[ 255] <= 6'h00;
      write_address_data_log_force[ 256] <= 6'h00;
      write_address_data_log_force[ 257] <= 6'h00;
      write_address_data_log_force[ 258] <= 6'h00;
      write_address_data_log_force[ 259] <= 6'h00;
      write_address_data_log_force[ 260] <= 6'h00;
      write_address_data_log_force[ 261] <= 6'h00;
      write_address_data_log_force[ 262] <= 6'h00;
      write_address_data_log_force[ 263] <= 6'h00;
      write_address_data_log_force[ 264] <= 6'h00;
      write_address_data_log_force[ 265] <= 6'h00;
      write_address_data_log_force[ 266] <= 6'h00;
      write_address_data_log_force[ 267] <= 6'h00;
      write_address_data_log_force[ 268] <= 6'h00;
      write_address_data_log_force[ 269] <= 6'h00;
      write_address_data_log_force[ 270] <= 6'h00;
      write_address_data_log_force[ 271] <= 6'h00;
      write_address_data_log_force[ 272] <= 6'h00;
      write_address_data_log_force[ 273] <= 6'h00;
      write_address_data_log_force[ 274] <= 6'h00;
      write_address_data_log_force[ 275] <= 6'h00;
      write_address_data_log_force[ 276] <= 6'h00;
      write_address_data_log_force[ 277] <= 6'h00;
      write_address_data_log_force[ 278] <= 6'h00;
      write_address_data_log_force[ 279] <= 6'h00;
      write_address_data_log_force[ 280] <= 6'h00;
      write_address_data_log_force[ 281] <= 6'h00;
      write_address_data_log_force[ 282] <= 6'h00;
      write_address_data_log_force[ 283] <= 6'h00;
      write_address_data_log_force[ 284] <= 6'h00;
      write_address_data_log_force[ 285] <= 6'h00;
      write_address_data_log_force[ 286] <= 6'h00;
      write_address_data_log_force[ 287] <= 6'h00;
      write_address_data_log_force[ 288] <= 6'h00;
      write_address_data_log_force[ 289] <= 6'h00;
      write_address_data_log_force[ 290] <= 6'h00;
      write_address_data_log_force[ 291] <= 6'h00;
      write_address_data_log_force[ 292] <= 6'h00;
      write_address_data_log_force[ 293] <= 6'h00;
      write_address_data_log_force[ 294] <= 6'h00;
      write_address_data_log_force[ 295] <= 6'h00;
      write_address_data_log_force[ 296] <= 6'h00;
      write_address_data_log_force[ 297] <= 6'h00;
      write_address_data_log_force[ 298] <= 6'h00;
      write_address_data_log_force[ 299] <= 6'h00;
      write_address_data_log_force[ 300] <= 6'h00;
      write_address_data_log_force[ 301] <= 6'h00;
      write_address_data_log_force[ 302] <= 6'h00;
      write_address_data_log_force[ 303] <= 6'h00;
      write_address_data_log_force[ 304] <= 6'h00;
      write_address_data_log_force[ 305] <= 6'h00;
      write_address_data_log_force[ 306] <= 6'h00;
      write_address_data_log_force[ 307] <= 6'h00;
      write_address_data_log_force[ 308] <= 6'h00;
      write_address_data_log_force[ 309] <= 6'h00;
      write_address_data_log_force[ 310] <= 6'h00;
      write_address_data_log_force[ 311] <= 6'h00;
      write_address_data_log_force[ 312] <= 6'h00;
      write_address_data_log_force[ 313] <= 6'h00;
      write_address_data_log_force[ 314] <= 6'h00;
      write_address_data_log_force[ 315] <= 6'h00;
      write_address_data_log_force[ 316] <= 6'h00;
      write_address_data_log_force[ 317] <= 6'h00;
      write_address_data_log_force[ 318] <= 6'h00;
      write_address_data_log_force[ 319] <= 6'h00;
      write_address_data_log_force[ 320] <= 6'h00;
      write_address_data_log_force[ 321] <= 6'h00;
      write_address_data_log_force[ 322] <= 6'h00;
      write_address_data_log_force[ 323] <= 6'h00;
      write_address_data_log_force[ 324] <= 6'h00;
      write_address_data_log_force[ 325] <= 6'h00;
      write_address_data_log_force[ 326] <= 6'h00;
      write_address_data_log_force[ 327] <= 6'h00;
      write_address_data_log_force[ 328] <= 6'h00;
      write_address_data_log_force[ 329] <= 6'h00;
      write_address_data_log_force[ 330] <= 6'h00;
      write_address_data_log_force[ 331] <= 6'h00;
      write_address_data_log_force[ 332] <= 6'h00;
      write_address_data_log_force[ 333] <= 6'h00;
      write_address_data_log_force[ 334] <= 6'h00;
      write_address_data_log_force[ 335] <= 6'h00;
      write_address_data_log_force[ 336] <= 6'h00;
      write_address_data_log_force[ 337] <= 6'h00;
      write_address_data_log_force[ 338] <= 6'h00;
      write_address_data_log_force[ 339] <= 6'h00;
      write_address_data_log_force[ 340] <= 6'h00;
      write_address_data_log_force[ 341] <= 6'h00;
      write_address_data_log_force[ 342] <= 6'h00;
      write_address_data_log_force[ 343] <= 6'h00;
      write_address_data_log_force[ 344] <= 6'h00;
      write_address_data_log_force[ 345] <= 6'h00;
      write_address_data_log_force[ 346] <= 6'h00;
      write_address_data_log_force[ 347] <= 6'h00;
      write_address_data_log_force[ 348] <= 6'h00;
      write_address_data_log_force[ 349] <= 6'h00;
      write_address_data_log_force[ 350] <= 6'h00;
      write_address_data_log_force[ 351] <= 6'h00;
      write_address_data_log_force[ 352] <= 6'h00;
      write_address_data_log_force[ 353] <= 6'h00;
      write_address_data_log_force[ 354] <= 6'h00;
      write_address_data_log_force[ 355] <= 6'h00;
      write_address_data_log_force[ 356] <= 6'h00;
      write_address_data_log_force[ 357] <= 6'h00;
      write_address_data_log_force[ 358] <= 6'h00;
      write_address_data_log_force[ 359] <= 6'h00;
      write_address_data_log_force[ 360] <= 6'h00;
      write_address_data_log_force[ 361] <= 6'h00;
      write_address_data_log_force[ 362] <= 6'h00;
      write_address_data_log_force[ 363] <= 6'h00;
      write_address_data_log_force[ 364] <= 6'h00;
      write_address_data_log_force[ 365] <= 6'h00;
      write_address_data_log_force[ 366] <= 6'h00;
      write_address_data_log_force[ 367] <= 6'h00;
      write_address_data_log_force[ 368] <= 6'h00;
      write_address_data_log_force[ 369] <= 6'h00;
      write_address_data_log_force[ 370] <= 6'h00;
      write_address_data_log_force[ 371] <= 6'h00;
      write_address_data_log_force[ 372] <= 6'h00;
      write_address_data_log_force[ 373] <= 6'h00;
      write_address_data_log_force[ 374] <= 6'h00;
      write_address_data_log_force[ 375] <= 6'h00;
      write_address_data_log_force[ 376] <= 6'h00;
      write_address_data_log_force[ 377] <= 6'h00;
      write_address_data_log_force[ 378] <= 6'h00;
      write_address_data_log_force[ 379] <= 6'h00;
      write_address_data_log_force[ 380] <= 6'h00;
      write_address_data_log_force[ 381] <= 6'h00;
      write_address_data_log_force[ 382] <= 6'h00;
      write_address_data_log_force[ 383] <= 6'h00;
      write_address_data_log_force[ 384] <= 6'h00;
      write_address_data_log_force[ 385] <= 6'h00;
      write_address_data_log_force[ 386] <= 6'h00;
      write_address_data_log_force[ 387] <= 6'h00;
      write_address_data_log_force[ 388] <= 6'h00;
      write_address_data_log_force[ 389] <= 6'h00;
      write_address_data_log_force[ 390] <= 6'h00;
      write_address_data_log_force[ 391] <= 6'h00;
      write_address_data_log_force[ 392] <= 6'h00;
      write_address_data_log_force[ 393] <= 6'h00;
      write_address_data_log_force[ 394] <= 6'h00;
      write_address_data_log_force[ 395] <= 6'h00;
      write_address_data_log_force[ 396] <= 6'h00;
      write_address_data_log_force[ 397] <= 6'h00;
      write_address_data_log_force[ 398] <= 6'h00;
      write_address_data_log_force[ 399] <= 6'h00;
      write_address_data_log_force[ 400] <= 6'h00;
      write_address_data_log_force[ 401] <= 6'h00;
      write_address_data_log_force[ 402] <= 6'h00;
      write_address_data_log_force[ 403] <= 6'h00;
      write_address_data_log_force[ 404] <= 6'h00;
      write_address_data_log_force[ 405] <= 6'h00;
      write_address_data_log_force[ 406] <= 6'h00;
      write_address_data_log_force[ 407] <= 6'h00;
      write_address_data_log_force[ 408] <= 6'h00;
      write_address_data_log_force[ 409] <= 6'h00;
      write_address_data_log_force[ 410] <= 6'h00;
      write_address_data_log_force[ 411] <= 6'h00;
      write_address_data_log_force[ 412] <= 6'h00;
      write_address_data_log_force[ 413] <= 6'h00;
      write_address_data_log_force[ 414] <= 6'h00;
      write_address_data_log_force[ 415] <= 6'h00;
      write_address_data_log_force[ 416] <= 6'h00;
      write_address_data_log_force[ 417] <= 6'h00;
      write_address_data_log_force[ 418] <= 6'h00;
      write_address_data_log_force[ 419] <= 6'h00;
      write_address_data_log_force[ 420] <= 6'h00;
      write_address_data_log_force[ 421] <= 6'h00;
      write_address_data_log_force[ 422] <= 6'h00;
      write_address_data_log_force[ 423] <= 6'h00;
      write_address_data_log_force[ 424] <= 6'h00;
      write_address_data_log_force[ 425] <= 6'h00;
      write_address_data_log_force[ 426] <= 6'h00;
      write_address_data_log_force[ 427] <= 6'h00;
      write_address_data_log_force[ 428] <= 6'h00;
      write_address_data_log_force[ 429] <= 6'h00;
      write_address_data_log_force[ 430] <= 6'h00;
      write_address_data_log_force[ 431] <= 6'h00;
      write_address_data_log_force[ 432] <= 6'h00;
      write_address_data_log_force[ 433] <= 6'h00;
      write_address_data_log_force[ 434] <= 6'h00;
      write_address_data_log_force[ 435] <= 6'h00;
      write_address_data_log_force[ 436] <= 6'h00;
      write_address_data_log_force[ 437] <= 6'h00;
      write_address_data_log_force[ 438] <= 6'h00;
      write_address_data_log_force[ 439] <= 6'h00;
      write_address_data_log_force[ 440] <= 6'h00;
      write_address_data_log_force[ 441] <= 6'h00;
      write_address_data_log_force[ 442] <= 6'h00;
      write_address_data_log_force[ 443] <= 6'h00;
      write_address_data_log_force[ 444] <= 6'h00;
      write_address_data_log_force[ 445] <= 6'h00;
      write_address_data_log_force[ 446] <= 6'h00;
      write_address_data_log_force[ 447] <= 6'h00;
      write_address_data_log_force[ 448] <= 6'h00;
      write_address_data_log_force[ 449] <= 6'h00;
      write_address_data_log_force[ 450] <= 6'h00;
      write_address_data_log_force[ 451] <= 6'h00;
      write_address_data_log_force[ 452] <= 6'h00;
      write_address_data_log_force[ 453] <= 6'h00;
      write_address_data_log_force[ 454] <= 6'h00;
      write_address_data_log_force[ 455] <= 6'h00;
      write_address_data_log_force[ 456] <= 6'h00;
      write_address_data_log_force[ 457] <= 6'h00;
      write_address_data_log_force[ 458] <= 6'h00;
      write_address_data_log_force[ 459] <= 6'h00;
      write_address_data_log_force[ 460] <= 6'h00;
      write_address_data_log_force[ 461] <= 6'h00;
      write_address_data_log_force[ 462] <= 6'h00;
      write_address_data_log_force[ 463] <= 6'h00;
      write_address_data_log_force[ 464] <= 6'h00;
      write_address_data_log_force[ 465] <= 6'h00;
      write_address_data_log_force[ 466] <= 6'h00;
      write_address_data_log_force[ 467] <= 6'h00;
      write_address_data_log_force[ 468] <= 6'h00;
      write_address_data_log_force[ 469] <= 6'h00;
      write_address_data_log_force[ 470] <= 6'h00;
      write_address_data_log_force[ 471] <= 6'h00;
      write_address_data_log_force[ 472] <= 6'h00;
      write_address_data_log_force[ 473] <= 6'h00;
      write_address_data_log_force[ 474] <= 6'h00;
      write_address_data_log_force[ 475] <= 6'h00;
      write_address_data_log_force[ 476] <= 6'h00;
      write_address_data_log_force[ 477] <= 6'h00;
      write_address_data_log_force[ 478] <= 6'h00;
      write_address_data_log_force[ 479] <= 6'h00;
      write_address_data_log_force[ 480] <= 6'h00;
      write_address_data_log_force[ 481] <= 6'h00;
      write_address_data_log_force[ 482] <= 6'h00;
      write_address_data_log_force[ 483] <= 6'h00;
      write_address_data_log_force[ 484] <= 6'h00;
      write_address_data_log_force[ 485] <= 6'h00;
      write_address_data_log_force[ 486] <= 6'h00;
      write_address_data_log_force[ 487] <= 6'h00;
      write_address_data_log_force[ 488] <= 6'h00;
      write_address_data_log_force[ 489] <= 6'h00;
      write_address_data_log_force[ 490] <= 6'h00;
      write_address_data_log_force[ 491] <= 6'h00;
      write_address_data_log_force[ 492] <= 6'h00;
      write_address_data_log_force[ 493] <= 6'h00;
      write_address_data_log_force[ 494] <= 6'h00;
      write_address_data_log_force[ 495] <= 6'h00;
      write_address_data_log_force[ 496] <= 6'h00;
      write_address_data_log_force[ 497] <= 6'h00;
      write_address_data_log_force[ 498] <= 6'h00;
      write_address_data_log_force[ 499] <= 6'h00;
      write_address_data_log_force[ 500] <= 6'h00;
      write_address_data_log_force[ 501] <= 6'h00;
      write_address_data_log_force[ 502] <= 6'h00;
      write_address_data_log_force[ 503] <= 6'h00;
      write_address_data_log_force[ 504] <= 6'h00;
      write_address_data_log_force[ 505] <= 6'h00;
      write_address_data_log_force[ 506] <= 6'h00;
      write_address_data_log_force[ 507] <= 6'h00;
      write_address_data_log_force[ 508] <= 6'h00;
      write_address_data_log_force[ 509] <= 6'h00;
      write_address_data_log_force[ 510] <= 6'h00;
      write_address_data_log_force[ 511] <= 6'h00;
      write_address_data_log_force[ 512] <= 6'h00;
      write_address_data_log_force[ 513] <= 6'h00;
      write_address_data_log_force[ 514] <= 6'h00;
      write_address_data_log_force[ 515] <= 6'h00;
      write_address_data_log_force[ 516] <= 6'h00;
      write_address_data_log_force[ 517] <= 6'h00;
      write_address_data_log_force[ 518] <= 6'h00;
      write_address_data_log_force[ 519] <= 6'h00;
      write_address_data_log_force[ 520] <= 6'h00;
      write_address_data_log_force[ 521] <= 6'h00;
      write_address_data_log_force[ 522] <= 6'h00;
      write_address_data_log_force[ 523] <= 6'h00;
      write_address_data_log_force[ 524] <= 6'h00;
      write_address_data_log_force[ 525] <= 6'h00;
      write_address_data_log_force[ 526] <= 6'h00;
      write_address_data_log_force[ 527] <= 6'h00;
      write_address_data_log_force[ 528] <= 6'h00;
      write_address_data_log_force[ 529] <= 6'h00;
      write_address_data_log_force[ 530] <= 6'h00;
      write_address_data_log_force[ 531] <= 6'h00;
      write_address_data_log_force[ 532] <= 6'h00;
      write_address_data_log_force[ 533] <= 6'h00;
      write_address_data_log_force[ 534] <= 6'h00;
      write_address_data_log_force[ 535] <= 6'h00;
      write_address_data_log_force[ 536] <= 6'h00;
      write_address_data_log_force[ 537] <= 6'h00;
      write_address_data_log_force[ 538] <= 6'h00;
      write_address_data_log_force[ 539] <= 6'h00;
      write_address_data_log_force[ 540] <= 6'h00;
      write_address_data_log_force[ 541] <= 6'h00;
      write_address_data_log_force[ 542] <= 6'h00;
      write_address_data_log_force[ 543] <= 6'h00;
      write_address_data_log_force[ 544] <= 6'h00;
      write_address_data_log_force[ 545] <= 6'h00;
      write_address_data_log_force[ 546] <= 6'h00;
      write_address_data_log_force[ 547] <= 6'h00;
      write_address_data_log_force[ 548] <= 6'h00;
      write_address_data_log_force[ 549] <= 6'h00;
      write_address_data_log_force[ 550] <= 6'h00;
      write_address_data_log_force[ 551] <= 6'h00;
      write_address_data_log_force[ 552] <= 6'h00;
      write_address_data_log_force[ 553] <= 6'h00;
      write_address_data_log_force[ 554] <= 6'h00;
      write_address_data_log_force[ 555] <= 6'h00;
      write_address_data_log_force[ 556] <= 6'h00;
      write_address_data_log_force[ 557] <= 6'h00;
      write_address_data_log_force[ 558] <= 6'h00;
      write_address_data_log_force[ 559] <= 6'h00;
      write_address_data_log_force[ 560] <= 6'h00;
      write_address_data_log_force[ 561] <= 6'h00;
      write_address_data_log_force[ 562] <= 6'h00;
      write_address_data_log_force[ 563] <= 6'h00;
      write_address_data_log_force[ 564] <= 6'h00;
      write_address_data_log_force[ 565] <= 6'h00;
      write_address_data_log_force[ 566] <= 6'h00;
      write_address_data_log_force[ 567] <= 6'h00;
      write_address_data_log_force[ 568] <= 6'h00;
      write_address_data_log_force[ 569] <= 6'h00;
      write_address_data_log_force[ 570] <= 6'h00;
      write_address_data_log_force[ 571] <= 6'h00;
      write_address_data_log_force[ 572] <= 6'h00;
      write_address_data_log_force[ 573] <= 6'h00;
      write_address_data_log_force[ 574] <= 6'h00;
      write_address_data_log_force[ 575] <= 6'h00;
      write_address_data_log_force[ 576] <= 6'h00;
      write_address_data_log_force[ 577] <= 6'h00;
      write_address_data_log_force[ 578] <= 6'h00;
      write_address_data_log_force[ 579] <= 6'h00;
      write_address_data_log_force[ 580] <= 6'h00;
      write_address_data_log_force[ 581] <= 6'h00;
      write_address_data_log_force[ 582] <= 6'h00;
      write_address_data_log_force[ 583] <= 6'h00;
      write_address_data_log_force[ 584] <= 6'h00;
      write_address_data_log_force[ 585] <= 6'h00;
      write_address_data_log_force[ 586] <= 6'h00;
      write_address_data_log_force[ 587] <= 6'h00;
      write_address_data_log_force[ 588] <= 6'h00;
      write_address_data_log_force[ 589] <= 6'h00;
      write_address_data_log_force[ 590] <= 6'h00;
      write_address_data_log_force[ 591] <= 6'h00;
      write_address_data_log_force[ 592] <= 6'h00;
      write_address_data_log_force[ 593] <= 6'h00;
      write_address_data_log_force[ 594] <= 6'h00;
      write_address_data_log_force[ 595] <= 6'h00;
      write_address_data_log_force[ 596] <= 6'h00;
      write_address_data_log_force[ 597] <= 6'h00;
      write_address_data_log_force[ 598] <= 6'h00;
      write_address_data_log_force[ 599] <= 6'h00;
      write_address_data_log_force[ 600] <= 6'h00;
      write_address_data_log_force[ 601] <= 6'h00;
      write_address_data_log_force[ 602] <= 6'h00;
      write_address_data_log_force[ 603] <= 6'h00;
      write_address_data_log_force[ 604] <= 6'h00;
      write_address_data_log_force[ 605] <= 6'h00;
      write_address_data_log_force[ 606] <= 6'h00;
      write_address_data_log_force[ 607] <= 6'h00;
      write_address_data_log_force[ 608] <= 6'h00;
      write_address_data_log_force[ 609] <= 6'h00;
      write_address_data_log_force[ 610] <= 6'h00;
      write_address_data_log_force[ 611] <= 6'h00;
      write_address_data_log_force[ 612] <= 6'h00;
      write_address_data_log_force[ 613] <= 6'h00;
      write_address_data_log_force[ 614] <= 6'h00;
      write_address_data_log_force[ 615] <= 6'h00;
      write_address_data_log_force[ 616] <= 6'h00;
      write_address_data_log_force[ 617] <= 6'h00;
      write_address_data_log_force[ 618] <= 6'h00;
      write_address_data_log_force[ 619] <= 6'h00;
      write_address_data_log_force[ 620] <= 6'h00;
      write_address_data_log_force[ 621] <= 6'h00;
      write_address_data_log_force[ 622] <= 6'h00;
      write_address_data_log_force[ 623] <= 6'h00;
      write_address_data_log_force[ 624] <= 6'h00;
      write_address_data_log_force[ 625] <= 6'h00;
      write_address_data_log_force[ 626] <= 6'h00;
      write_address_data_log_force[ 627] <= 6'h00;
      write_address_data_log_force[ 628] <= 6'h00;
      write_address_data_log_force[ 629] <= 6'h00;
      write_address_data_log_force[ 630] <= 6'h00;
      write_address_data_log_force[ 631] <= 6'h00;
      write_address_data_log_force[ 632] <= 6'h00;
      write_address_data_log_force[ 633] <= 6'h00;
      write_address_data_log_force[ 634] <= 6'h00;
      write_address_data_log_force[ 635] <= 6'h00;
      write_address_data_log_force[ 636] <= 6'h00;
      write_address_data_log_force[ 637] <= 6'h00;
      write_address_data_log_force[ 638] <= 6'h00;
      write_address_data_log_force[ 639] <= 6'h00;
      write_address_data_log_force[ 640] <= 6'h00;
      write_address_data_log_force[ 641] <= 6'h00;
      write_address_data_log_force[ 642] <= 6'h00;
      write_address_data_log_force[ 643] <= 6'h00;
      write_address_data_log_force[ 644] <= 6'h00;
      write_address_data_log_force[ 645] <= 6'h00;
      write_address_data_log_force[ 646] <= 6'h00;
      write_address_data_log_force[ 647] <= 6'h00;
      write_address_data_log_force[ 648] <= 6'h00;
      write_address_data_log_force[ 649] <= 6'h00;
      write_address_data_log_force[ 650] <= 6'h00;
      write_address_data_log_force[ 651] <= 6'h00;
      write_address_data_log_force[ 652] <= 6'h00;
      write_address_data_log_force[ 653] <= 6'h00;
      write_address_data_log_force[ 654] <= 6'h00;
      write_address_data_log_force[ 655] <= 6'h00;
      write_address_data_log_force[ 656] <= 6'h00;
      write_address_data_log_force[ 657] <= 6'h00;
      write_address_data_log_force[ 658] <= 6'h00;
      write_address_data_log_force[ 659] <= 6'h00;
      write_address_data_log_force[ 660] <= 6'h00;
      write_address_data_log_force[ 661] <= 6'h00;
      write_address_data_log_force[ 662] <= 6'h00;
      write_address_data_log_force[ 663] <= 6'h00;
      write_address_data_log_force[ 664] <= 6'h00;
      write_address_data_log_force[ 665] <= 6'h00;
      write_address_data_log_force[ 666] <= 6'h00;
      write_address_data_log_force[ 667] <= 6'h00;
      write_address_data_log_force[ 668] <= 6'h00;
      write_address_data_log_force[ 669] <= 6'h00;
      write_address_data_log_force[ 670] <= 6'h00;
      write_address_data_log_force[ 671] <= 6'h00;
      write_address_data_log_force[ 672] <= 6'h00;
      write_address_data_log_force[ 673] <= 6'h00;
      write_address_data_log_force[ 674] <= 6'h00;
      write_address_data_log_force[ 675] <= 6'h00;
      write_address_data_log_force[ 676] <= 6'h00;
      write_address_data_log_force[ 677] <= 6'h00;
      write_address_data_log_force[ 678] <= 6'h00;
      write_address_data_log_force[ 679] <= 6'h00;
      write_address_data_log_force[ 680] <= 6'h00;
      write_address_data_log_force[ 681] <= 6'h00;
      write_address_data_log_force[ 682] <= 6'h00;
      write_address_data_log_force[ 683] <= 6'h00;
      write_address_data_log_force[ 684] <= 6'h00;
      write_address_data_log_force[ 685] <= 6'h00;
      write_address_data_log_force[ 686] <= 6'h00;
      write_address_data_log_force[ 687] <= 6'h00;
      write_address_data_log_force[ 688] <= 6'h00;
      write_address_data_log_force[ 689] <= 6'h00;
      write_address_data_log_force[ 690] <= 6'h00;
      write_address_data_log_force[ 691] <= 6'h00;
      write_address_data_log_force[ 692] <= 6'h00;
      write_address_data_log_force[ 693] <= 6'h00;
      write_address_data_log_force[ 694] <= 6'h00;
      write_address_data_log_force[ 695] <= 6'h00;
      write_address_data_log_force[ 696] <= 6'h00;
      write_address_data_log_force[ 697] <= 6'h00;
      write_address_data_log_force[ 698] <= 6'h00;
      write_address_data_log_force[ 699] <= 6'h00;
      write_address_data_log_force[ 700] <= 6'h00;
      write_address_data_log_force[ 701] <= 6'h00;
      write_address_data_log_force[ 702] <= 6'h00;
      write_address_data_log_force[ 703] <= 6'h00;
      write_address_data_log_force[ 704] <= 6'h00;
      write_address_data_log_force[ 705] <= 6'h00;
      write_address_data_log_force[ 706] <= 6'h00;
      write_address_data_log_force[ 707] <= 6'h00;
      write_address_data_log_force[ 708] <= 6'h00;
      write_address_data_log_force[ 709] <= 6'h00;
      write_address_data_log_force[ 710] <= 6'h00;
      write_address_data_log_force[ 711] <= 6'h00;
      write_address_data_log_force[ 712] <= 6'h00;
      write_address_data_log_force[ 713] <= 6'h00;
      write_address_data_log_force[ 714] <= 6'h00;
      write_address_data_log_force[ 715] <= 6'h00;
      write_address_data_log_force[ 716] <= 6'h00;
      write_address_data_log_force[ 717] <= 6'h00;
      write_address_data_log_force[ 718] <= 6'h00;
      write_address_data_log_force[ 719] <= 6'h00;
      write_address_data_log_force[ 720] <= 6'h00;
      write_address_data_log_force[ 721] <= 6'h00;
      write_address_data_log_force[ 722] <= 6'h00;
      write_address_data_log_force[ 723] <= 6'h00;
      write_address_data_log_force[ 724] <= 6'h00;
      write_address_data_log_force[ 725] <= 6'h00;
      write_address_data_log_force[ 726] <= 6'h00;
      write_address_data_log_force[ 727] <= 6'h00;
      write_address_data_log_force[ 728] <= 6'h00;
      write_address_data_log_force[ 729] <= 6'h00;
      write_address_data_log_force[ 730] <= 6'h00;
      write_address_data_log_force[ 731] <= 6'h00;
      write_address_data_log_force[ 732] <= 6'h00;
      write_address_data_log_force[ 733] <= 6'h00;
      write_address_data_log_force[ 734] <= 6'h00;
      write_address_data_log_force[ 735] <= 6'h00;
      write_address_data_log_force[ 736] <= 6'h00;
      write_address_data_log_force[ 737] <= 6'h00;
      write_address_data_log_force[ 738] <= 6'h00;
      write_address_data_log_force[ 739] <= 6'h00;
      write_address_data_log_force[ 740] <= 6'h00;
      write_address_data_log_force[ 741] <= 6'h00;
      write_address_data_log_force[ 742] <= 6'h00;
      write_address_data_log_force[ 743] <= 6'h00;
      write_address_data_log_force[ 744] <= 6'h00;
      write_address_data_log_force[ 745] <= 6'h00;
      write_address_data_log_force[ 746] <= 6'h00;
      write_address_data_log_force[ 747] <= 6'h00;
      write_address_data_log_force[ 748] <= 6'h00;
      write_address_data_log_force[ 749] <= 6'h00;
      write_address_data_log_force[ 750] <= 6'h00;
      write_address_data_log_force[ 751] <= 6'h00;
      write_address_data_log_force[ 752] <= 6'h00;
      write_address_data_log_force[ 753] <= 6'h00;
      write_address_data_log_force[ 754] <= 6'h00;
      write_address_data_log_force[ 755] <= 6'h00;
      write_address_data_log_force[ 756] <= 6'h00;
      write_address_data_log_force[ 757] <= 6'h00;
      write_address_data_log_force[ 758] <= 6'h00;
      write_address_data_log_force[ 759] <= 6'h00;
      write_address_data_log_force[ 760] <= 6'h00;
      write_address_data_log_force[ 761] <= 6'h00;
      write_address_data_log_force[ 762] <= 6'h00;
      write_address_data_log_force[ 763] <= 6'h00;
      write_address_data_log_force[ 764] <= 6'h00;
      write_address_data_log_force[ 765] <= 6'h00;
      write_address_data_log_force[ 766] <= 6'h00;
      write_address_data_log_force[ 767] <= 6'h00;
      write_address_data_log_force[ 768] <= 6'h00;
      write_address_data_log_force[ 769] <= 6'h00;
      write_address_data_log_force[ 770] <= 6'h00;
      write_address_data_log_force[ 771] <= 6'h00;
      write_address_data_log_force[ 772] <= 6'h00;
      write_address_data_log_force[ 773] <= 6'h00;
      write_address_data_log_force[ 774] <= 6'h00;
      write_address_data_log_force[ 775] <= 6'h00;
      write_address_data_log_force[ 776] <= 6'h00;
      write_address_data_log_force[ 777] <= 6'h00;
      write_address_data_log_force[ 778] <= 6'h00;
      write_address_data_log_force[ 779] <= 6'h00;
      write_address_data_log_force[ 780] <= 6'h00;
      write_address_data_log_force[ 781] <= 6'h00;
      write_address_data_log_force[ 782] <= 6'h00;
      write_address_data_log_force[ 783] <= 6'h00;
      write_address_data_log_force[ 784] <= 6'h00;
      write_address_data_log_force[ 785] <= 6'h00;
      write_address_data_log_force[ 786] <= 6'h00;
      write_address_data_log_force[ 787] <= 6'h00;
      write_address_data_log_force[ 788] <= 6'h00;
      write_address_data_log_force[ 789] <= 6'h00;
      write_address_data_log_force[ 790] <= 6'h00;
      write_address_data_log_force[ 791] <= 6'h00;
      write_address_data_log_force[ 792] <= 6'h00;
      write_address_data_log_force[ 793] <= 6'h00;
      write_address_data_log_force[ 794] <= 6'h00;
      write_address_data_log_force[ 795] <= 6'h00;
      write_address_data_log_force[ 796] <= 6'h00;
      write_address_data_log_force[ 797] <= 6'h00;
      write_address_data_log_force[ 798] <= 6'h00;
      write_address_data_log_force[ 799] <= 6'h00;
      write_address_data_log_force[ 800] <= 6'h00;
      write_address_data_log_force[ 801] <= 6'h00;
      write_address_data_log_force[ 802] <= 6'h00;
      write_address_data_log_force[ 803] <= 6'h00;
      write_address_data_log_force[ 804] <= 6'h00;
      write_address_data_log_force[ 805] <= 6'h00;
      write_address_data_log_force[ 806] <= 6'h00;
      write_address_data_log_force[ 807] <= 6'h00;
      write_address_data_log_force[ 808] <= 6'h00;
      write_address_data_log_force[ 809] <= 6'h00;
      write_address_data_log_force[ 810] <= 6'h00;
      write_address_data_log_force[ 811] <= 6'h00;
      write_address_data_log_force[ 812] <= 6'h00;
      write_address_data_log_force[ 813] <= 6'h00;
      write_address_data_log_force[ 814] <= 6'h00;
      write_address_data_log_force[ 815] <= 6'h00;
      write_address_data_log_force[ 816] <= 6'h00;
      write_address_data_log_force[ 817] <= 6'h00;
      write_address_data_log_force[ 818] <= 6'h00;
      write_address_data_log_force[ 819] <= 6'h00;
      write_address_data_log_force[ 820] <= 6'h00;
      write_address_data_log_force[ 821] <= 6'h00;
      write_address_data_log_force[ 822] <= 6'h00;
      write_address_data_log_force[ 823] <= 6'h00;
      write_address_data_log_force[ 824] <= 6'h00;
      write_address_data_log_force[ 825] <= 6'h00;
      write_address_data_log_force[ 826] <= 6'h00;
      write_address_data_log_force[ 827] <= 6'h00;
      write_address_data_log_force[ 828] <= 6'h00;
      write_address_data_log_force[ 829] <= 6'h00;
      write_address_data_log_force[ 830] <= 6'h00;
      write_address_data_log_force[ 831] <= 6'h00;
      write_address_data_log_force[ 832] <= 6'h00;
      write_address_data_log_force[ 833] <= 6'h00;
      write_address_data_log_force[ 834] <= 6'h00;
      write_address_data_log_force[ 835] <= 6'h00;
      write_address_data_log_force[ 836] <= 6'h00;
      write_address_data_log_force[ 837] <= 6'h00;
      write_address_data_log_force[ 838] <= 6'h00;
      write_address_data_log_force[ 839] <= 6'h00;
      write_address_data_log_force[ 840] <= 6'h00;
      write_address_data_log_force[ 841] <= 6'h00;
      write_address_data_log_force[ 842] <= 6'h00;
      write_address_data_log_force[ 843] <= 6'h00;
      write_address_data_log_force[ 844] <= 6'h00;
      write_address_data_log_force[ 845] <= 6'h00;
      write_address_data_log_force[ 846] <= 6'h00;
      write_address_data_log_force[ 847] <= 6'h00;
      write_address_data_log_force[ 848] <= 6'h00;
      write_address_data_log_force[ 849] <= 6'h00;
      write_address_data_log_force[ 850] <= 6'h00;
      write_address_data_log_force[ 851] <= 6'h00;
      write_address_data_log_force[ 852] <= 6'h00;
      write_address_data_log_force[ 853] <= 6'h00;
      write_address_data_log_force[ 854] <= 6'h00;
      write_address_data_log_force[ 855] <= 6'h00;
      write_address_data_log_force[ 856] <= 6'h00;
      write_address_data_log_force[ 857] <= 6'h00;
      write_address_data_log_force[ 858] <= 6'h00;
      write_address_data_log_force[ 859] <= 6'h00;
      write_address_data_log_force[ 860] <= 6'h00;
      write_address_data_log_force[ 861] <= 6'h00;
      write_address_data_log_force[ 862] <= 6'h00;
      write_address_data_log_force[ 863] <= 6'h00;
      write_address_data_log_force[ 864] <= 6'h00;
      write_address_data_log_force[ 865] <= 6'h00;
      write_address_data_log_force[ 866] <= 6'h00;
      write_address_data_log_force[ 867] <= 6'h00;
      write_address_data_log_force[ 868] <= 6'h00;
      write_address_data_log_force[ 869] <= 6'h00;
      write_address_data_log_force[ 870] <= 6'h00;
      write_address_data_log_force[ 871] <= 6'h00;
      write_address_data_log_force[ 872] <= 6'h00;
      write_address_data_log_force[ 873] <= 6'h00;
      write_address_data_log_force[ 874] <= 6'h00;
      write_address_data_log_force[ 875] <= 6'h00;
      write_address_data_log_force[ 876] <= 6'h00;
      write_address_data_log_force[ 877] <= 6'h00;
      write_address_data_log_force[ 878] <= 6'h00;
      write_address_data_log_force[ 879] <= 6'h00;
      write_address_data_log_force[ 880] <= 6'h00;
      write_address_data_log_force[ 881] <= 6'h00;
      write_address_data_log_force[ 882] <= 6'h00;
      write_address_data_log_force[ 883] <= 6'h00;
      write_address_data_log_force[ 884] <= 6'h00;
      write_address_data_log_force[ 885] <= 6'h00;
      write_address_data_log_force[ 886] <= 6'h00;
      write_address_data_log_force[ 887] <= 6'h00;
      write_address_data_log_force[ 888] <= 6'h00;
      write_address_data_log_force[ 889] <= 6'h00;
      write_address_data_log_force[ 890] <= 6'h00;
      write_address_data_log_force[ 891] <= 6'h00;
      write_address_data_log_force[ 892] <= 6'h00;
      write_address_data_log_force[ 893] <= 6'h00;
      write_address_data_log_force[ 894] <= 6'h00;
      write_address_data_log_force[ 895] <= 6'h00;
      write_address_data_log_force[ 896] <= 6'h00;
      write_address_data_log_force[ 897] <= 6'h00;
      write_address_data_log_force[ 898] <= 6'h00;
      write_address_data_log_force[ 899] <= 6'h00;
      write_address_data_log_force[ 900] <= 6'h00;
      write_address_data_log_force[ 901] <= 6'h00;
      write_address_data_log_force[ 902] <= 6'h00;
      write_address_data_log_force[ 903] <= 6'h00;
      write_address_data_log_force[ 904] <= 6'h00;
      write_address_data_log_force[ 905] <= 6'h00;
      write_address_data_log_force[ 906] <= 6'h00;
      write_address_data_log_force[ 907] <= 6'h00;
      write_address_data_log_force[ 908] <= 6'h00;
      write_address_data_log_force[ 909] <= 6'h00;
      write_address_data_log_force[ 910] <= 6'h00;
      write_address_data_log_force[ 911] <= 6'h00;
      write_address_data_log_force[ 912] <= 6'h00;
      write_address_data_log_force[ 913] <= 6'h00;
      write_address_data_log_force[ 914] <= 6'h00;
      write_address_data_log_force[ 915] <= 6'h00;
      write_address_data_log_force[ 916] <= 6'h00;
      write_address_data_log_force[ 917] <= 6'h00;
      write_address_data_log_force[ 918] <= 6'h00;
      write_address_data_log_force[ 919] <= 6'h00;
      write_address_data_log_force[ 920] <= 6'h00;
      write_address_data_log_force[ 921] <= 6'h00;
      write_address_data_log_force[ 922] <= 6'h00;
      write_address_data_log_force[ 923] <= 6'h00;
      write_address_data_log_force[ 924] <= 6'h00;
      write_address_data_log_force[ 925] <= 6'h00;
      write_address_data_log_force[ 926] <= 6'h00;
      write_address_data_log_force[ 927] <= 6'h00;
      write_address_data_log_force[ 928] <= 6'h00;
      write_address_data_log_force[ 929] <= 6'h00;
      write_address_data_log_force[ 930] <= 6'h00;
      write_address_data_log_force[ 931] <= 6'h00;
      write_address_data_log_force[ 932] <= 6'h00;
      write_address_data_log_force[ 933] <= 6'h00;
      write_address_data_log_force[ 934] <= 6'h00;
      write_address_data_log_force[ 935] <= 6'h00;
      write_address_data_log_force[ 936] <= 6'h00;
      write_address_data_log_force[ 937] <= 6'h00;
      write_address_data_log_force[ 938] <= 6'h00;
      write_address_data_log_force[ 939] <= 6'h00;
      write_address_data_log_force[ 940] <= 6'h00;
      write_address_data_log_force[ 941] <= 6'h00;
      write_address_data_log_force[ 942] <= 6'h00;
      write_address_data_log_force[ 943] <= 6'h00;
      write_address_data_log_force[ 944] <= 6'h00;
      write_address_data_log_force[ 945] <= 6'h00;
      write_address_data_log_force[ 946] <= 6'h00;
      write_address_data_log_force[ 947] <= 6'h00;
      write_address_data_log_force[ 948] <= 6'h00;
      write_address_data_log_force[ 949] <= 6'h00;
      write_address_data_log_force[ 950] <= 6'h00;
      write_address_data_log_force[ 951] <= 6'h00;
      write_address_data_log_force[ 952] <= 6'h00;
      write_address_data_log_force[ 953] <= 6'h00;
      write_address_data_log_force[ 954] <= 6'h00;
      write_address_data_log_force[ 955] <= 6'h00;
      write_address_data_log_force[ 956] <= 6'h00;
      write_address_data_log_force[ 957] <= 6'h00;
      write_address_data_log_force[ 958] <= 6'h00;
      write_address_data_log_force[ 959] <= 6'h00;
      write_address_data_log_force[ 960] <= 6'h00;
      write_address_data_log_force[ 961] <= 6'h00;
      write_address_data_log_force[ 962] <= 6'h00;
      write_address_data_log_force[ 963] <= 6'h00;
      write_address_data_log_force[ 964] <= 6'h00;
      write_address_data_log_force[ 965] <= 6'h00;
      write_address_data_log_force[ 966] <= 6'h00;
      write_address_data_log_force[ 967] <= 6'h00;
      write_address_data_log_force[ 968] <= 6'h00;
      write_address_data_log_force[ 969] <= 6'h00;
      write_address_data_log_force[ 970] <= 6'h00;
      write_address_data_log_force[ 971] <= 6'h00;
      write_address_data_log_force[ 972] <= 6'h00;
      write_address_data_log_force[ 973] <= 6'h00;
      write_address_data_log_force[ 974] <= 6'h00;
      write_address_data_log_force[ 975] <= 6'h00;
      write_address_data_log_force[ 976] <= 6'h00;
      write_address_data_log_force[ 977] <= 6'h00;
      write_address_data_log_force[ 978] <= 6'h00;
      write_address_data_log_force[ 979] <= 6'h00;
      write_address_data_log_force[ 980] <= 6'h00;
      write_address_data_log_force[ 981] <= 6'h00;
      write_address_data_log_force[ 982] <= 6'h00;
      write_address_data_log_force[ 983] <= 6'h00;
      write_address_data_log_force[ 984] <= 6'h00;
      write_address_data_log_force[ 985] <= 6'h00;
      write_address_data_log_force[ 986] <= 6'h00;
      write_address_data_log_force[ 987] <= 6'h00;
      write_address_data_log_force[ 988] <= 6'h00;
      write_address_data_log_force[ 989] <= 6'h00;
      write_address_data_log_force[ 990] <= 6'h00;
      write_address_data_log_force[ 991] <= 6'h00;
      write_address_data_log_force[ 992] <= 6'h00;
      write_address_data_log_force[ 993] <= 6'h00;
      write_address_data_log_force[ 994] <= 6'h00;
      write_address_data_log_force[ 995] <= 6'h00;
      write_address_data_log_force[ 996] <= 6'h00;
      write_address_data_log_force[ 997] <= 6'h00;
      write_address_data_log_force[ 998] <= 6'h00;
      write_address_data_log_force[ 999] <= 6'h00;
      write_address_data_log_force[1000] <= 6'h00;
      write_address_data_log_force[1001] <= 6'h00;
      write_address_data_log_force[1002] <= 6'h00;
      write_address_data_log_force[1003] <= 6'h00;
      write_address_data_log_force[1004] <= 6'h00;
      write_address_data_log_force[1005] <= 6'h00;
      write_address_data_log_force[1006] <= 6'h00;
      write_address_data_log_force[1007] <= 6'h00;
      write_address_data_log_force[1008] <= 6'h00;
      write_address_data_log_force[1009] <= 6'h00;
      write_address_data_log_force[1010] <= 6'h00;
      write_address_data_log_force[1011] <= 6'h00;
      write_address_data_log_force[1012] <= 6'h00;
      write_address_data_log_force[1013] <= 6'h00;
      write_address_data_log_force[1014] <= 6'h00;
      write_address_data_log_force[1015] <= 6'h00;
      write_address_data_log_force[1016] <= 6'h00;
      write_address_data_log_force[1017] <= 6'h00;
      write_address_data_log_force[1018] <= 6'h00;
      write_address_data_log_force[1019] <= 6'h00;
      write_address_data_log_force[1020] <= 6'h00;
      write_address_data_log_force[1021] <= 6'h00;
      write_address_data_log_force[1022] <= 6'h00;
      write_address_data_log_force[1023] <= 6'h00;
      write_address_data_log_force[1024] <= 6'h00;
      write_address_data_log_force[1025] <= 6'h00;
      write_address_data_log_force[1026] <= 6'h00;
      write_address_data_log_force[1027] <= 6'h00;
      write_address_data_log_force[1028] <= 6'h00;
      write_address_data_log_force[1029] <= 6'h00;
      write_address_data_log_force[1030] <= 6'h00;
      write_address_data_log_force[1031] <= 6'h00;
      write_address_data_log_force[1032] <= 6'h00;
      write_address_data_log_force[1033] <= 6'h00;
      write_address_data_log_force[1034] <= 6'h00;
      write_address_data_log_force[1035] <= 6'h00;
      write_address_data_log_force[1036] <= 6'h00;
      write_address_data_log_force[1037] <= 6'h00;
      write_address_data_log_force[1038] <= 6'h00;
      write_address_data_log_force[1039] <= 6'h00;
      write_address_data_log_force[1040] <= 6'h00;
      write_address_data_log_force[1041] <= 6'h00;
      write_address_data_log_force[1042] <= 6'h00;
      write_address_data_log_force[1043] <= 6'h00;
      write_address_data_log_force[1044] <= 6'h00;
      write_address_data_log_force[1045] <= 6'h00;
      write_address_data_log_force[1046] <= 6'h00;
      write_address_data_log_force[1047] <= 6'h00;
      write_address_data_log_force[1048] <= 6'h00;
      write_address_data_log_force[1049] <= 6'h00;
      write_address_data_log_force[1050] <= 6'h00;
      write_address_data_log_force[1051] <= 6'h00;
      write_address_data_log_force[1052] <= 6'h00;
      write_address_data_log_force[1053] <= 6'h00;
      write_address_data_log_force[1054] <= 6'h00;
      write_address_data_log_force[1055] <= 6'h00;
      write_address_data_log_force[1056] <= 6'h00;
      write_address_data_log_force[1057] <= 6'h00;
      write_address_data_log_force[1058] <= 6'h00;
      write_address_data_log_force[1059] <= 6'h00;
      write_address_data_log_force[1060] <= 6'h00;
      write_address_data_log_force[1061] <= 6'h00;
      write_address_data_log_force[1062] <= 6'h00;
      write_address_data_log_force[1063] <= 6'h00;
      write_address_data_log_force[1064] <= 6'h00;
      write_address_data_log_force[1065] <= 6'h00;
      write_address_data_log_force[1066] <= 6'h00;
      write_address_data_log_force[1067] <= 6'h00;
      write_address_data_log_force[1068] <= 6'h00;
      write_address_data_log_force[1069] <= 6'h00;
      write_address_data_log_force[1070] <= 6'h00;
      write_address_data_log_force[1071] <= 6'h00;
      write_address_data_log_force[1072] <= 6'h00;
      write_address_data_log_force[1073] <= 6'h00;
      write_address_data_log_force[1074] <= 6'h00;
      write_address_data_log_force[1075] <= 6'h00;
      write_address_data_log_force[1076] <= 6'h00;
      write_address_data_log_force[1077] <= 6'h00;
      write_address_data_log_force[1078] <= 6'h00;
      write_address_data_log_force[1079] <= 6'h00;
      write_address_data_log_force[1080] <= 6'h00;
      write_address_data_log_force[1081] <= 6'h00;
      write_address_data_log_force[1082] <= 6'h00;
      write_address_data_log_force[1083] <= 6'h00;
      write_address_data_log_force[1084] <= 6'h00;
      write_address_data_log_force[1085] <= 6'h00;
      write_address_data_log_force[1086] <= 6'h00;
      write_address_data_log_force[1087] <= 6'h00;
      write_address_data_log_force[1088] <= 6'h00;
      write_address_data_log_force[1089] <= 6'h00;
      write_address_data_log_force[1090] <= 6'h00;
      write_address_data_log_force[1091] <= 6'h00;
      write_address_data_log_force[1092] <= 6'h00;
      write_address_data_log_force[1093] <= 6'h00;
      write_address_data_log_force[1094] <= 6'h00;
      write_address_data_log_force[1095] <= 6'h00;
      write_address_data_log_force[1096] <= 6'h00;
      write_address_data_log_force[1097] <= 6'h00;
      write_address_data_log_force[1098] <= 6'h00;
      write_address_data_log_force[1099] <= 6'h00;
      write_address_data_log_force[1100] <= 6'h00;
      write_address_data_log_force[1101] <= 6'h00;
      write_address_data_log_force[1102] <= 6'h00;
      write_address_data_log_force[1103] <= 6'h00;
      write_address_data_log_force[1104] <= 6'h00;
      write_address_data_log_force[1105] <= 6'h00;
      write_address_data_log_force[1106] <= 6'h00;
      write_address_data_log_force[1107] <= 6'h00;
      write_address_data_log_force[1108] <= 6'h00;
      write_address_data_log_force[1109] <= 6'h00;
      write_address_data_log_force[1110] <= 6'h00;
      write_address_data_log_force[1111] <= 6'h00;
      write_address_data_log_force[1112] <= 6'h00;
      write_address_data_log_force[1113] <= 6'h00;
      write_address_data_log_force[1114] <= 6'h00;
      write_address_data_log_force[1115] <= 6'h00;
      write_address_data_log_force[1116] <= 6'h00;
      write_address_data_log_force[1117] <= 6'h00;
      write_address_data_log_force[1118] <= 6'h00;
      write_address_data_log_force[1119] <= 6'h00;
      write_address_data_log_force[1120] <= 6'h00;
      write_address_data_log_force[1121] <= 6'h00;
      write_address_data_log_force[1122] <= 6'h00;
      write_address_data_log_force[1123] <= 6'h00;
      write_address_data_log_force[1124] <= 6'h00;
      write_address_data_log_force[1125] <= 6'h00;
      write_address_data_log_force[1126] <= 6'h00;
      write_address_data_log_force[1127] <= 6'h00;
      write_address_data_log_force[1128] <= 6'h00;
      write_address_data_log_force[1129] <= 6'h00;
      write_address_data_log_force[1130] <= 6'h00;
      write_address_data_log_force[1131] <= 6'h00;
      write_address_data_log_force[1132] <= 6'h00;
      write_address_data_log_force[1133] <= 6'h00;
      write_address_data_log_force[1134] <= 6'h00;
      write_address_data_log_force[1135] <= 6'h00;
      write_address_data_log_force[1136] <= 6'h00;
      write_address_data_log_force[1137] <= 6'h00;
      write_address_data_log_force[1138] <= 6'h00;
      write_address_data_log_force[1139] <= 6'h00;
      write_address_data_log_force[1140] <= 6'h00;
      write_address_data_log_force[1141] <= 6'h00;
      write_address_data_log_force[1142] <= 6'h00;
      write_address_data_log_force[1143] <= 6'h00;
      write_address_data_log_force[1144] <= 6'h00;
      write_address_data_log_force[1145] <= 6'h00;
      write_address_data_log_force[1146] <= 6'h00;
      write_address_data_log_force[1147] <= 6'h00;
      write_address_data_log_force[1148] <= 6'h00;
      write_address_data_log_force[1149] <= 6'h00;
      write_address_data_log_force[1150] <= 6'h00;
      write_address_data_log_force[1151] <= 6'h00;
      write_address_data_log_force[1152] <= 6'h00;
      write_address_data_log_force[1153] <= 6'h00;
      write_address_data_log_force[1154] <= 6'h00;
      write_address_data_log_force[1155] <= 6'h00;
      write_address_data_log_force[1156] <= 6'h00;
      write_address_data_log_force[1157] <= 6'h00;
      write_address_data_log_force[1158] <= 6'h00;
      write_address_data_log_force[1159] <= 6'h00;
      write_address_data_log_force[1160] <= 6'h00;
      write_address_data_log_force[1161] <= 6'h00;
      write_address_data_log_force[1162] <= 6'h00;
      write_address_data_log_force[1163] <= 6'h00;
      write_address_data_log_force[1164] <= 6'h00;
      write_address_data_log_force[1165] <= 6'h00;
      write_address_data_log_force[1166] <= 6'h00;
      write_address_data_log_force[1167] <= 6'h00;
      write_address_data_log_force[1168] <= 6'h00;
      write_address_data_log_force[1169] <= 6'h00;
      write_address_data_log_force[1170] <= 6'h00;
      write_address_data_log_force[1171] <= 6'h00;
      write_address_data_log_force[1172] <= 6'h00;
      write_address_data_log_force[1173] <= 6'h00;
      write_address_data_log_force[1174] <= 6'h00;
      write_address_data_log_force[1175] <= 6'h00;
      write_address_data_log_force[1176] <= 6'h00;
      write_address_data_log_force[1177] <= 6'h00;
      write_address_data_log_force[1178] <= 6'h00;
      write_address_data_log_force[1179] <= 6'h00;
      write_address_data_log_force[1180] <= 6'h00;
      write_address_data_log_force[1181] <= 6'h00;
      write_address_data_log_force[1182] <= 6'h00;
      write_address_data_log_force[1183] <= 6'h00;
      write_address_data_log_force[1184] <= 6'h00;
      write_address_data_log_force[1185] <= 6'h00;
      write_address_data_log_force[1186] <= 6'h00;
      write_address_data_log_force[1187] <= 6'h00;
      write_address_data_log_force[1188] <= 6'h00;
      write_address_data_log_force[1189] <= 6'h00;
      write_address_data_log_force[1190] <= 6'h00;
      write_address_data_log_force[1191] <= 6'h00;
      write_address_data_log_force[1192] <= 6'h00;
      write_address_data_log_force[1193] <= 6'h00;
      write_address_data_log_force[1194] <= 6'h00;
      write_address_data_log_force[1195] <= 6'h00;
      write_address_data_log_force[1196] <= 6'h00;
      write_address_data_log_force[1197] <= 6'h00;
      write_address_data_log_force[1198] <= 6'h00;
      write_address_data_log_force[1199] <= 6'h00;
      write_address_data_log_force[1200] <= 6'h00;
      write_address_data_log_force[1201] <= 6'h00;
      write_address_data_log_force[1202] <= 6'h00;
      write_address_data_log_force[1203] <= 6'h00;
      write_address_data_log_force[1204] <= 6'h00;
      write_address_data_log_force[1205] <= 6'h00;
      write_address_data_log_force[1206] <= 6'h00;
      write_address_data_log_force[1207] <= 6'h00;
      write_address_data_log_force[1208] <= 6'h00;
      write_address_data_log_force[1209] <= 6'h00;
      write_address_data_log_force[1210] <= 6'h00;
      write_address_data_log_force[1211] <= 6'h00;
      write_address_data_log_force[1212] <= 6'h00;
      write_address_data_log_force[1213] <= 6'h00;
      write_address_data_log_force[1214] <= 6'h00;
      write_address_data_log_force[1215] <= 6'h00;
      write_address_data_log_force[1216] <= 6'h00;
      write_address_data_log_force[1217] <= 6'h00;
      write_address_data_log_force[1218] <= 6'h00;
      write_address_data_log_force[1219] <= 6'h00;
      write_address_data_log_force[1220] <= 6'h00;
      write_address_data_log_force[1221] <= 6'h00;
      write_address_data_log_force[1222] <= 6'h00;
      write_address_data_log_force[1223] <= 6'h00;
      write_address_data_log_force[1224] <= 6'h00;
      write_address_data_log_force[1225] <= 6'h00;
      write_address_data_log_force[1226] <= 6'h00;
      write_address_data_log_force[1227] <= 6'h00;
      write_address_data_log_force[1228] <= 6'h00;
      write_address_data_log_force[1229] <= 6'h00;
      write_address_data_log_force[1230] <= 6'h00;
      write_address_data_log_force[1231] <= 6'h00;
      write_address_data_log_force[1232] <= 6'h00;
      write_address_data_log_force[1233] <= 6'h00;
      write_address_data_log_force[1234] <= 6'h00;
      write_address_data_log_force[1235] <= 6'h00;
      write_address_data_log_force[1236] <= 6'h00;
      write_address_data_log_force[1237] <= 6'h00;
      write_address_data_log_force[1238] <= 6'h00;
      write_address_data_log_force[1239] <= 6'h00;
      write_address_data_log_force[1240] <= 6'h00;
      write_address_data_log_force[1241] <= 6'h00;
      write_address_data_log_force[1242] <= 6'h00;
      write_address_data_log_force[1243] <= 6'h00;
      write_address_data_log_force[1244] <= 6'h00;
      write_address_data_log_force[1245] <= 6'h00;
      write_address_data_log_force[1246] <= 6'h00;
      write_address_data_log_force[1247] <= 6'h00;
      write_address_data_log_force[1248] <= 6'h00;
      write_address_data_log_force[1249] <= 6'h00;
      write_address_data_log_force[1250] <= 6'h00;
      write_address_data_log_force[1251] <= 6'h00;
      write_address_data_log_force[1252] <= 6'h00;
      write_address_data_log_force[1253] <= 6'h00;
      write_address_data_log_force[1254] <= 6'h00;
      write_address_data_log_force[1255] <= 6'h00;
      write_address_data_log_force[1256] <= 6'h00;
      write_address_data_log_force[1257] <= 6'h00;
      write_address_data_log_force[1258] <= 6'h00;
      write_address_data_log_force[1259] <= 6'h00;
      write_address_data_log_force[1260] <= 6'h00;
      write_address_data_log_force[1261] <= 6'h00;
      write_address_data_log_force[1262] <= 6'h00;
      write_address_data_log_force[1263] <= 6'h00;
      write_address_data_log_force[1264] <= 6'h00;
      write_address_data_log_force[1265] <= 6'h00;
      write_address_data_log_force[1266] <= 6'h00;
      write_address_data_log_force[1267] <= 6'h00;
      write_address_data_log_force[1268] <= 6'h00;
      write_address_data_log_force[1269] <= 6'h00;
      write_address_data_log_force[1270] <= 6'h00;
      write_address_data_log_force[1271] <= 6'h00;
      write_address_data_log_force[1272] <= 6'h00;
      write_address_data_log_force[1273] <= 6'h00;
      write_address_data_log_force[1274] <= 6'h00;
      write_address_data_log_force[1275] <= 6'h00;
      write_address_data_log_force[1276] <= 6'h00;
      write_address_data_log_force[1277] <= 6'h00;
      write_address_data_log_force[1278] <= 6'h00;
      write_address_data_log_force[1279] <= 6'h00;
      write_address_data_log_force[1280] <= 6'h00;
      write_address_data_log_force[1281] <= 6'h00;
      write_address_data_log_force[1282] <= 6'h00;
      write_address_data_log_force[1283] <= 6'h00;
      write_address_data_log_force[1284] <= 6'h00;
      write_address_data_log_force[1285] <= 6'h00;
      write_address_data_log_force[1286] <= 6'h00;
      write_address_data_log_force[1287] <= 6'h00;
      write_address_data_log_force[1288] <= 6'h00;
      write_address_data_log_force[1289] <= 6'h00;
      write_address_data_log_force[1290] <= 6'h00;
      write_address_data_log_force[1291] <= 6'h00;
      write_address_data_log_force[1292] <= 6'h00;
      write_address_data_log_force[1293] <= 6'h00;
      write_address_data_log_force[1294] <= 6'h00;
      write_address_data_log_force[1295] <= 6'h00;
      write_address_data_log_force[1296] <= 6'h00;
      write_address_data_log_force[1297] <= 6'h00;
      write_address_data_log_force[1298] <= 6'h00;
      write_address_data_log_force[1299] <= 6'h00;
      write_address_data_log_force[1300] <= 6'h00;
      write_address_data_log_force[1301] <= 6'h00;
      write_address_data_log_force[1302] <= 6'h00;
      write_address_data_log_force[1303] <= 6'h00;
      write_address_data_log_force[1304] <= 6'h00;
      write_address_data_log_force[1305] <= 6'h00;
      write_address_data_log_force[1306] <= 6'h00;
      write_address_data_log_force[1307] <= 6'h00;
      write_address_data_log_force[1308] <= 6'h00;
      write_address_data_log_force[1309] <= 6'h00;
      write_address_data_log_force[1310] <= 6'h00;
      write_address_data_log_force[1311] <= 6'h00;
      write_address_data_log_force[1312] <= 6'h00;
      write_address_data_log_force[1313] <= 6'h00;
      write_address_data_log_force[1314] <= 6'h00;
      write_address_data_log_force[1315] <= 6'h00;
      write_address_data_log_force[1316] <= 6'h00;
      write_address_data_log_force[1317] <= 6'h00;
      write_address_data_log_force[1318] <= 6'h00;
      write_address_data_log_force[1319] <= 6'h00;
      write_address_data_log_force[1320] <= 6'h00;
      write_address_data_log_force[1321] <= 6'h00;
      write_address_data_log_force[1322] <= 6'h00;
      write_address_data_log_force[1323] <= 6'h00;
      write_address_data_log_force[1324] <= 6'h00;
      write_address_data_log_force[1325] <= 6'h00;
      write_address_data_log_force[1326] <= 6'h00;
      write_address_data_log_force[1327] <= 6'h00;
      write_address_data_log_force[1328] <= 6'h00;
      write_address_data_log_force[1329] <= 6'h00;
      write_address_data_log_force[1330] <= 6'h00;
      write_address_data_log_force[1331] <= 6'h00;
      write_address_data_log_force[1332] <= 6'h00;
      write_address_data_log_force[1333] <= 6'h00;
      write_address_data_log_force[1334] <= 6'h00;
      write_address_data_log_force[1335] <= 6'h00;
      write_address_data_log_force[1336] <= 6'h00;
      write_address_data_log_force[1337] <= 6'h00;
      write_address_data_log_force[1338] <= 6'h00;
      write_address_data_log_force[1339] <= 6'h00;
      write_address_data_log_force[1340] <= 6'h00;
      write_address_data_log_force[1341] <= 6'h00;
      write_address_data_log_force[1342] <= 6'h00;
      write_address_data_log_force[1343] <= 6'h00;
      write_address_data_log_force[1344] <= 6'h00;
      write_address_data_log_force[1345] <= 6'h00;
      write_address_data_log_force[1346] <= 6'h00;
      write_address_data_log_force[1347] <= 6'h00;
      write_address_data_log_force[1348] <= 6'h00;
      write_address_data_log_force[1349] <= 6'h00;
      write_address_data_log_force[1350] <= 6'h00;
      write_address_data_log_force[1351] <= 6'h00;
      write_address_data_log_force[1352] <= 6'h00;
      write_address_data_log_force[1353] <= 6'h00;
      write_address_data_log_force[1354] <= 6'h00;
      write_address_data_log_force[1355] <= 6'h00;
      write_address_data_log_force[1356] <= 6'h00;
      write_address_data_log_force[1357] <= 6'h00;
      write_address_data_log_force[1358] <= 6'h00;
      write_address_data_log_force[1359] <= 6'h00;
      write_address_data_log_force[1360] <= 6'h00;
      write_address_data_log_force[1361] <= 6'h00;
      write_address_data_log_force[1362] <= 6'h00;
      write_address_data_log_force[1363] <= 6'h00;
      write_address_data_log_force[1364] <= 6'h00;
      write_address_data_log_force[1365] <= 6'h00;
      write_address_data_log_force[1366] <= 6'h00;
      write_address_data_log_force[1367] <= 6'h00;
      write_address_data_log_force[1368] <= 6'h00;
      write_address_data_log_force[1369] <= 6'h00;
      write_address_data_log_force[1370] <= 6'h00;
      write_address_data_log_force[1371] <= 6'h00;
      write_address_data_log_force[1372] <= 6'h00;
      write_address_data_log_force[1373] <= 6'h00;
      write_address_data_log_force[1374] <= 6'h00;
      write_address_data_log_force[1375] <= 6'h00;
      write_address_data_log_force[1376] <= 6'h00;
      write_address_data_log_force[1377] <= 6'h00;
      write_address_data_log_force[1378] <= 6'h00;
      write_address_data_log_force[1379] <= 6'h00;
      write_address_data_log_force[1380] <= 6'h00;
      write_address_data_log_force[1381] <= 6'h00;
      write_address_data_log_force[1382] <= 6'h00;
      write_address_data_log_force[1383] <= 6'h00;
      write_address_data_log_force[1384] <= 6'h00;
      write_address_data_log_force[1385] <= 6'h00;
      write_address_data_log_force[1386] <= 6'h00;
      write_address_data_log_force[1387] <= 6'h00;
      write_address_data_log_force[1388] <= 6'h00;
      write_address_data_log_force[1389] <= 6'h00;
      write_address_data_log_force[1390] <= 6'h00;
      write_address_data_log_force[1391] <= 6'h00;
      write_address_data_log_force[1392] <= 6'h00;
      write_address_data_log_force[1393] <= 6'h00;
      write_address_data_log_force[1394] <= 6'h00;
      write_address_data_log_force[1395] <= 6'h00;
      write_address_data_log_force[1396] <= 6'h00;
      write_address_data_log_force[1397] <= 6'h00;
      write_address_data_log_force[1398] <= 6'h00;
      write_address_data_log_force[1399] <= 6'h00;
      write_address_data_log_force[1400] <= 6'h00;
      write_address_data_log_force[1401] <= 6'h00;
      write_address_data_log_force[1402] <= 6'h00;
      write_address_data_log_force[1403] <= 6'h00;
      write_address_data_log_force[1404] <= 6'h00;
      write_address_data_log_force[1405] <= 6'h00;
      write_address_data_log_force[1406] <= 6'h00;
      write_address_data_log_force[1407] <= 6'h00;
      write_address_data_log_force[1408] <= 6'h00;
      write_address_data_log_force[1409] <= 6'h00;
      write_address_data_log_force[1410] <= 6'h00;
      write_address_data_log_force[1411] <= 6'h00;
      write_address_data_log_force[1412] <= 6'h00;
      write_address_data_log_force[1413] <= 6'h00;
      write_address_data_log_force[1414] <= 6'h00;
      write_address_data_log_force[1415] <= 6'h00;
      write_address_data_log_force[1416] <= 6'h00;
      write_address_data_log_force[1417] <= 6'h00;
      write_address_data_log_force[1418] <= 6'h00;
      write_address_data_log_force[1419] <= 6'h00;
      write_address_data_log_force[1420] <= 6'h00;
      write_address_data_log_force[1421] <= 6'h00;
      write_address_data_log_force[1422] <= 6'h00;
      write_address_data_log_force[1423] <= 6'h00;
      write_address_data_log_force[1424] <= 6'h00;
      write_address_data_log_force[1425] <= 6'h00;
      write_address_data_log_force[1426] <= 6'h00;
      write_address_data_log_force[1427] <= 6'h00;
      write_address_data_log_force[1428] <= 6'h00;
      write_address_data_log_force[1429] <= 6'h00;
      write_address_data_log_force[1430] <= 6'h00;
      write_address_data_log_force[1431] <= 6'h00;
      write_address_data_log_force[1432] <= 6'h00;
      write_address_data_log_force[1433] <= 6'h00;
      write_address_data_log_force[1434] <= 6'h00;
      write_address_data_log_force[1435] <= 6'h00;
      write_address_data_log_force[1436] <= 6'h00;
      write_address_data_log_force[1437] <= 6'h00;
      write_address_data_log_force[1438] <= 6'h00;
      write_address_data_log_force[1439] <= 6'h00;
      write_address_data_log_force[1440] <= 6'h00;
      write_address_data_log_force[1441] <= 6'h00;
      write_address_data_log_force[1442] <= 6'h00;
      write_address_data_log_force[1443] <= 6'h00;
      write_address_data_log_force[1444] <= 6'h00;
      write_address_data_log_force[1445] <= 6'h00;
      write_address_data_log_force[1446] <= 6'h00;
      write_address_data_log_force[1447] <= 6'h00;
      write_address_data_log_force[1448] <= 6'h00;
      write_address_data_log_force[1449] <= 6'h00;
      write_address_data_log_force[1450] <= 6'h00;
      write_address_data_log_force[1451] <= 6'h00;
      write_address_data_log_force[1452] <= 6'h00;
      write_address_data_log_force[1453] <= 6'h00;
      write_address_data_log_force[1454] <= 6'h00;
      write_address_data_log_force[1455] <= 6'h00;
      write_address_data_log_force[1456] <= 6'h00;
      write_address_data_log_force[1457] <= 6'h00;
      write_address_data_log_force[1458] <= 6'h00;
      write_address_data_log_force[1459] <= 6'h00;
      write_address_data_log_force[1460] <= 6'h00;
      write_address_data_log_force[1461] <= 6'h00;
      write_address_data_log_force[1462] <= 6'h00;
      write_address_data_log_force[1463] <= 6'h00;
      write_address_data_log_force[1464] <= 6'h00;
      write_address_data_log_force[1465] <= 6'h00;
      write_address_data_log_force[1466] <= 6'h00;
      write_address_data_log_force[1467] <= 6'h00;
      write_address_data_log_force[1468] <= 6'h00;
      write_address_data_log_force[1469] <= 6'h00;
      write_address_data_log_force[1470] <= 6'h00;
      write_address_data_log_force[1471] <= 6'h00;
      write_address_data_log_force[1472] <= 6'h00;
      write_address_data_log_force[1473] <= 6'h00;
      write_address_data_log_force[1474] <= 6'h00;
      write_address_data_log_force[1475] <= 6'h00;
      write_address_data_log_force[1476] <= 6'h00;
      write_address_data_log_force[1477] <= 6'h00;
      write_address_data_log_force[1478] <= 6'h00;
      write_address_data_log_force[1479] <= 6'h00;
      write_address_data_log_force[1480] <= 6'h00;
      write_address_data_log_force[1481] <= 6'h00;
      write_address_data_log_force[1482] <= 6'h00;
      write_address_data_log_force[1483] <= 6'h00;
      write_address_data_log_force[1484] <= 6'h00;
      write_address_data_log_force[1485] <= 6'h00;
      write_address_data_log_force[1486] <= 6'h00;
      write_address_data_log_force[1487] <= 6'h00;
      write_address_data_log_force[1488] <= 6'h00;
      write_address_data_log_force[1489] <= 6'h00;
      write_address_data_log_force[1490] <= 6'h00;
      write_address_data_log_force[1491] <= 6'h00;
      write_address_data_log_force[1492] <= 6'h00;
      write_address_data_log_force[1493] <= 6'h00;
      write_address_data_log_force[1494] <= 6'h00;
      write_address_data_log_force[1495] <= 6'h00;
      write_address_data_log_force[1496] <= 6'h00;
      write_address_data_log_force[1497] <= 6'h00;
      write_address_data_log_force[1498] <= 6'h00;
      write_address_data_log_force[1499] <= 6'h00;
      write_address_data_log_force[1500] <= 6'h00;
      write_address_data_log_force[1501] <= 6'h00;
      write_address_data_log_force[1502] <= 6'h00;
      write_address_data_log_force[1503] <= 6'h00;
      write_address_data_log_force[1504] <= 6'h00;
      write_address_data_log_force[1505] <= 6'h00;
      write_address_data_log_force[1506] <= 6'h00;
      write_address_data_log_force[1507] <= 6'h00;
      write_address_data_log_force[1508] <= 6'h00;
      write_address_data_log_force[1509] <= 6'h00;
      write_address_data_log_force[1510] <= 6'h00;
      write_address_data_log_force[1511] <= 6'h00;
      write_address_data_log_force[1512] <= 6'h00;
      write_address_data_log_force[1513] <= 6'h00;
      write_address_data_log_force[1514] <= 6'h00;
      write_address_data_log_force[1515] <= 6'h00;
      write_address_data_log_force[1516] <= 6'h00;
      write_address_data_log_force[1517] <= 6'h00;
      write_address_data_log_force[1518] <= 6'h00;
      write_address_data_log_force[1519] <= 6'h00;
      write_address_data_log_force[1520] <= 6'h00;
      write_address_data_log_force[1521] <= 6'h00;
      write_address_data_log_force[1522] <= 6'h00;
      write_address_data_log_force[1523] <= 6'h00;
      write_address_data_log_force[1524] <= 6'h00;
      write_address_data_log_force[1525] <= 6'h00;
      write_address_data_log_force[1526] <= 6'h00;
      write_address_data_log_force[1527] <= 6'h00;
      write_address_data_log_force[1528] <= 6'h00;
      write_address_data_log_force[1529] <= 6'h00;
      write_address_data_log_force[1530] <= 6'h00;
      write_address_data_log_force[1531] <= 6'h00;
      write_address_data_log_force[1532] <= 6'h00;
      write_address_data_log_force[1533] <= 6'h00;
      write_address_data_log_force[1534] <= 6'h00;
      write_address_data_log_force[1535] <= 6'h00;
      write_address_data_log_force[1536] <= 6'h00;
      write_address_data_log_force[1537] <= 6'h00;
      write_address_data_log_force[1538] <= 6'h00;
      write_address_data_log_force[1539] <= 6'h00;
      write_address_data_log_force[1540] <= 6'h00;
      write_address_data_log_force[1541] <= 6'h00;
      write_address_data_log_force[1542] <= 6'h00;
      write_address_data_log_force[1543] <= 6'h00;
      write_address_data_log_force[1544] <= 6'h00;
      write_address_data_log_force[1545] <= 6'h00;
      write_address_data_log_force[1546] <= 6'h00;
      write_address_data_log_force[1547] <= 6'h00;
      write_address_data_log_force[1548] <= 6'h00;
      write_address_data_log_force[1549] <= 6'h00;
      write_address_data_log_force[1550] <= 6'h00;
      write_address_data_log_force[1551] <= 6'h00;
      write_address_data_log_force[1552] <= 6'h00;
      write_address_data_log_force[1553] <= 6'h00;
      write_address_data_log_force[1554] <= 6'h00;
      write_address_data_log_force[1555] <= 6'h00;
      write_address_data_log_force[1556] <= 6'h00;
      write_address_data_log_force[1557] <= 6'h00;
      write_address_data_log_force[1558] <= 6'h00;
      write_address_data_log_force[1559] <= 6'h00;
      write_address_data_log_force[1560] <= 6'h00;
      write_address_data_log_force[1561] <= 6'h00;
      write_address_data_log_force[1562] <= 6'h00;
      write_address_data_log_force[1563] <= 6'h00;
      write_address_data_log_force[1564] <= 6'h00;
      write_address_data_log_force[1565] <= 6'h00;
      write_address_data_log_force[1566] <= 6'h00;
      write_address_data_log_force[1567] <= 6'h00;
      write_address_data_log_force[1568] <= 6'h00;
      write_address_data_log_force[1569] <= 6'h00;
      write_address_data_log_force[1570] <= 6'h00;
      write_address_data_log_force[1571] <= 6'h00;
      write_address_data_log_force[1572] <= 6'h00;
      write_address_data_log_force[1573] <= 6'h00;
      write_address_data_log_force[1574] <= 6'h00;
      write_address_data_log_force[1575] <= 6'h00;
      write_address_data_log_force[1576] <= 6'h00;
      write_address_data_log_force[1577] <= 6'h00;
      write_address_data_log_force[1578] <= 6'h00;
      write_address_data_log_force[1579] <= 6'h00;
      write_address_data_log_force[1580] <= 6'h00;
      write_address_data_log_force[1581] <= 6'h00;
      write_address_data_log_force[1582] <= 6'h00;
      write_address_data_log_force[1583] <= 6'h00;
      write_address_data_log_force[1584] <= 6'h00;
      write_address_data_log_force[1585] <= 6'h00;
      write_address_data_log_force[1586] <= 6'h00;
      write_address_data_log_force[1587] <= 6'h00;
      write_address_data_log_force[1588] <= 6'h00;
      write_address_data_log_force[1589] <= 6'h00;
      write_address_data_log_force[1590] <= 6'h00;
      write_address_data_log_force[1591] <= 6'h00;
      write_address_data_log_force[1592] <= 6'h00;
      write_address_data_log_force[1593] <= 6'h00;
      write_address_data_log_force[1594] <= 6'h00;
      write_address_data_log_force[1595] <= 6'h00;
      write_address_data_log_force[1596] <= 6'h00;
      write_address_data_log_force[1597] <= 6'h00;
      write_address_data_log_force[1598] <= 6'h00;
      write_address_data_log_force[1599] <= 6'h00;
      write_address_data_log_force[1600] <= 6'h00;
      write_address_data_log_force[1601] <= 6'h00;
      write_address_data_log_force[1602] <= 6'h00;
      write_address_data_log_force[1603] <= 6'h00;
      write_address_data_log_force[1604] <= 6'h00;
      write_address_data_log_force[1605] <= 6'h00;
      write_address_data_log_force[1606] <= 6'h00;
      write_address_data_log_force[1607] <= 6'h00;
      write_address_data_log_force[1608] <= 6'h00;
      write_address_data_log_force[1609] <= 6'h00;
      write_address_data_log_force[1610] <= 6'h00;
      write_address_data_log_force[1611] <= 6'h00;
      write_address_data_log_force[1612] <= 6'h00;
      write_address_data_log_force[1613] <= 6'h00;
      write_address_data_log_force[1614] <= 6'h00;
      write_address_data_log_force[1615] <= 6'h00;
      write_address_data_log_force[1616] <= 6'h00;
      write_address_data_log_force[1617] <= 6'h00;
      write_address_data_log_force[1618] <= 6'h00;
      write_address_data_log_force[1619] <= 6'h00;
      write_address_data_log_force[1620] <= 6'h00;
      write_address_data_log_force[1621] <= 6'h00;
      write_address_data_log_force[1622] <= 6'h00;
      write_address_data_log_force[1623] <= 6'h00;
      write_address_data_log_force[1624] <= 6'h00;
      write_address_data_log_force[1625] <= 6'h00;
      write_address_data_log_force[1626] <= 6'h00;
      write_address_data_log_force[1627] <= 6'h00;
      write_address_data_log_force[1628] <= 6'h00;
      write_address_data_log_force[1629] <= 6'h00;
      write_address_data_log_force[1630] <= 6'h00;
      write_address_data_log_force[1631] <= 6'h00;
      write_address_data_log_force[1632] <= 6'h00;
      write_address_data_log_force[1633] <= 6'h00;
      write_address_data_log_force[1634] <= 6'h00;
      write_address_data_log_force[1635] <= 6'h00;
      write_address_data_log_force[1636] <= 6'h00;
      write_address_data_log_force[1637] <= 6'h00;
      write_address_data_log_force[1638] <= 6'h00;
      write_address_data_log_force[1639] <= 6'h00;
      write_address_data_log_force[1640] <= 6'h00;
      write_address_data_log_force[1641] <= 6'h00;
      write_address_data_log_force[1642] <= 6'h00;
      write_address_data_log_force[1643] <= 6'h00;
      write_address_data_log_force[1644] <= 6'h00;
      write_address_data_log_force[1645] <= 6'h00;
      write_address_data_log_force[1646] <= 6'h00;
      write_address_data_log_force[1647] <= 6'h00;
      write_address_data_log_force[1648] <= 6'h00;
      write_address_data_log_force[1649] <= 6'h00;
      write_address_data_log_force[1650] <= 6'h00;
      write_address_data_log_force[1651] <= 6'h00;
      write_address_data_log_force[1652] <= 6'h00;
      write_address_data_log_force[1653] <= 6'h00;
      write_address_data_log_force[1654] <= 6'h00;
      write_address_data_log_force[1655] <= 6'h00;
      write_address_data_log_force[1656] <= 6'h00;
      write_address_data_log_force[1657] <= 6'h00;
      write_address_data_log_force[1658] <= 6'h00;
      write_address_data_log_force[1659] <= 6'h00;
      write_address_data_log_force[1660] <= 6'h00;
      write_address_data_log_force[1661] <= 6'h00;
      write_address_data_log_force[1662] <= 6'h00;
      write_address_data_log_force[1663] <= 6'h00;
      write_address_data_log_force[1664] <= 6'h00;
      write_address_data_log_force[1665] <= 6'h00;
      write_address_data_log_force[1666] <= 6'h00;
      write_address_data_log_force[1667] <= 6'h00;
      write_address_data_log_force[1668] <= 6'h00;
      write_address_data_log_force[1669] <= 6'h00;
      write_address_data_log_force[1670] <= 6'h00;
      write_address_data_log_force[1671] <= 6'h00;
      write_address_data_log_force[1672] <= 6'h00;
      write_address_data_log_force[1673] <= 6'h00;
      write_address_data_log_force[1674] <= 6'h00;
      write_address_data_log_force[1675] <= 6'h00;
      write_address_data_log_force[1676] <= 6'h00;
      write_address_data_log_force[1677] <= 6'h00;
      write_address_data_log_force[1678] <= 6'h00;
      write_address_data_log_force[1679] <= 6'h00;
      write_address_data_log_force[1680] <= 6'h00;
      write_address_data_log_force[1681] <= 6'h00;
      write_address_data_log_force[1682] <= 6'h00;
      write_address_data_log_force[1683] <= 6'h00;
      write_address_data_log_force[1684] <= 6'h00;
      write_address_data_log_force[1685] <= 6'h00;
      write_address_data_log_force[1686] <= 6'h00;
      write_address_data_log_force[1687] <= 6'h00;
      write_address_data_log_force[1688] <= 6'h00;
      write_address_data_log_force[1689] <= 6'h00;
      write_address_data_log_force[1690] <= 6'h00;
      write_address_data_log_force[1691] <= 6'h00;
      write_address_data_log_force[1692] <= 6'h00;
      write_address_data_log_force[1693] <= 6'h00;
      write_address_data_log_force[1694] <= 6'h00;
      write_address_data_log_force[1695] <= 6'h00;
      write_address_data_log_force[1696] <= 6'h00;
      write_address_data_log_force[1697] <= 6'h00;
      write_address_data_log_force[1698] <= 6'h00;
      write_address_data_log_force[1699] <= 6'h00;
      write_address_data_log_force[1700] <= 6'h00;
      write_address_data_log_force[1701] <= 6'h00;
      write_address_data_log_force[1702] <= 6'h00;
      write_address_data_log_force[1703] <= 6'h00;
      write_address_data_log_force[1704] <= 6'h00;
      write_address_data_log_force[1705] <= 6'h00;
      write_address_data_log_force[1706] <= 6'h00;
      write_address_data_log_force[1707] <= 6'h00;
      write_address_data_log_force[1708] <= 6'h00;
      write_address_data_log_force[1709] <= 6'h00;
      write_address_data_log_force[1710] <= 6'h00;
      write_address_data_log_force[1711] <= 6'h00;
      write_address_data_log_force[1712] <= 6'h00;
      write_address_data_log_force[1713] <= 6'h00;
      write_address_data_log_force[1714] <= 6'h00;
      write_address_data_log_force[1715] <= 6'h00;
      write_address_data_log_force[1716] <= 6'h00;
      write_address_data_log_force[1717] <= 6'h00;
      write_address_data_log_force[1718] <= 6'h00;
      write_address_data_log_force[1719] <= 6'h00;
      write_address_data_log_force[1720] <= 6'h00;
      write_address_data_log_force[1721] <= 6'h00;
      write_address_data_log_force[1722] <= 6'h00;
      write_address_data_log_force[1723] <= 6'h00;
      write_address_data_log_force[1724] <= 6'h00;
      write_address_data_log_force[1725] <= 6'h00;
      write_address_data_log_force[1726] <= 6'h00;
      write_address_data_log_force[1727] <= 6'h00;
      write_address_data_log_force[1728] <= 6'h00;
      write_address_data_log_force[1729] <= 6'h00;
      write_address_data_log_force[1730] <= 6'h00;
      write_address_data_log_force[1731] <= 6'h00;
      write_address_data_log_force[1732] <= 6'h00;
      write_address_data_log_force[1733] <= 6'h00;
      write_address_data_log_force[1734] <= 6'h00;
      write_address_data_log_force[1735] <= 6'h00;
      write_address_data_log_force[1736] <= 6'h00;
      write_address_data_log_force[1737] <= 6'h00;
      write_address_data_log_force[1738] <= 6'h00;
      write_address_data_log_force[1739] <= 6'h00;
      write_address_data_log_force[1740] <= 6'h00;
      write_address_data_log_force[1741] <= 6'h00;
      write_address_data_log_force[1742] <= 6'h00;
      write_address_data_log_force[1743] <= 6'h00;
      write_address_data_log_force[1744] <= 6'h00;
      write_address_data_log_force[1745] <= 6'h00;
      write_address_data_log_force[1746] <= 6'h00;
      write_address_data_log_force[1747] <= 6'h00;
      write_address_data_log_force[1748] <= 6'h00;
      write_address_data_log_force[1749] <= 6'h00;
      write_address_data_log_force[1750] <= 6'h00;
      write_address_data_log_force[1751] <= 6'h00;
      write_address_data_log_force[1752] <= 6'h00;
      write_address_data_log_force[1753] <= 6'h00;
      write_address_data_log_force[1754] <= 6'h00;
      write_address_data_log_force[1755] <= 6'h00;
      write_address_data_log_force[1756] <= 6'h00;
      write_address_data_log_force[1757] <= 6'h00;
      write_address_data_log_force[1758] <= 6'h00;
      write_address_data_log_force[1759] <= 6'h00;
      write_address_data_log_force[1760] <= 6'h00;
      write_address_data_log_force[1761] <= 6'h00;
      write_address_data_log_force[1762] <= 6'h00;
      write_address_data_log_force[1763] <= 6'h00;
      write_address_data_log_force[1764] <= 6'h00;
      write_address_data_log_force[1765] <= 6'h00;
      write_address_data_log_force[1766] <= 6'h00;
      write_address_data_log_force[1767] <= 6'h00;
      write_address_data_log_force[1768] <= 6'h00;
      write_address_data_log_force[1769] <= 6'h00;
      write_address_data_log_force[1770] <= 6'h00;
      write_address_data_log_force[1771] <= 6'h00;
      write_address_data_log_force[1772] <= 6'h00;
      write_address_data_log_force[1773] <= 6'h00;
      write_address_data_log_force[1774] <= 6'h00;
      write_address_data_log_force[1775] <= 6'h00;
      write_address_data_log_force[1776] <= 6'h00;
      write_address_data_log_force[1777] <= 6'h00;
      write_address_data_log_force[1778] <= 6'h00;
      write_address_data_log_force[1779] <= 6'h00;
      write_address_data_log_force[1780] <= 6'h00;
      write_address_data_log_force[1781] <= 6'h00;
      write_address_data_log_force[1782] <= 6'h00;
      write_address_data_log_force[1783] <= 6'h00;
      write_address_data_log_force[1784] <= 6'h00;
      write_address_data_log_force[1785] <= 6'h00;
      write_address_data_log_force[1786] <= 6'h00;
      write_address_data_log_force[1787] <= 6'h00;
      write_address_data_log_force[1788] <= 6'h00;
      write_address_data_log_force[1789] <= 6'h00;
      write_address_data_log_force[1790] <= 6'h00;
      write_address_data_log_force[1791] <= 6'h00;
      write_address_data_log_force[1792] <= 6'h00;
      write_address_data_log_force[1793] <= 6'h00;
      write_address_data_log_force[1794] <= 6'h00;
      write_address_data_log_force[1795] <= 6'h00;
      write_address_data_log_force[1796] <= 6'h00;
      write_address_data_log_force[1797] <= 6'h00;
      write_address_data_log_force[1798] <= 6'h00;
      write_address_data_log_force[1799] <= 6'h00;
      write_address_data_log_force[1800] <= 6'h00;
      write_address_data_log_force[1801] <= 6'h00;
      write_address_data_log_force[1802] <= 6'h00;
      write_address_data_log_force[1803] <= 6'h00;
      write_address_data_log_force[1804] <= 6'h00;
      write_address_data_log_force[1805] <= 6'h00;
      write_address_data_log_force[1806] <= 6'h00;
      write_address_data_log_force[1807] <= 6'h00;
      write_address_data_log_force[1808] <= 6'h00;
      write_address_data_log_force[1809] <= 6'h00;
      write_address_data_log_force[1810] <= 6'h00;
      write_address_data_log_force[1811] <= 6'h00;
      write_address_data_log_force[1812] <= 6'h00;
      write_address_data_log_force[1813] <= 6'h00;
      write_address_data_log_force[1814] <= 6'h00;
      write_address_data_log_force[1815] <= 6'h00;
      write_address_data_log_force[1816] <= 6'h00;
      write_address_data_log_force[1817] <= 6'h00;
      write_address_data_log_force[1818] <= 6'h00;
      write_address_data_log_force[1819] <= 6'h00;
      write_address_data_log_force[1820] <= 6'h00;
      write_address_data_log_force[1821] <= 6'h00;
      write_address_data_log_force[1822] <= 6'h00;
      write_address_data_log_force[1823] <= 6'h00;
      write_address_data_log_force[1824] <= 6'h00;
      write_address_data_log_force[1825] <= 6'h00;
      write_address_data_log_force[1826] <= 6'h00;
      write_address_data_log_force[1827] <= 6'h00;
      write_address_data_log_force[1828] <= 6'h00;
      write_address_data_log_force[1829] <= 6'h00;
      write_address_data_log_force[1830] <= 6'h00;
      write_address_data_log_force[1831] <= 6'h00;
      write_address_data_log_force[1832] <= 6'h00;
      write_address_data_log_force[1833] <= 6'h00;
      write_address_data_log_force[1834] <= 6'h00;
      write_address_data_log_force[1835] <= 6'h00;
      write_address_data_log_force[1836] <= 6'h00;
      write_address_data_log_force[1837] <= 6'h00;
      write_address_data_log_force[1838] <= 6'h00;
      write_address_data_log_force[1839] <= 6'h00;
      write_address_data_log_force[1840] <= 6'h00;
      write_address_data_log_force[1841] <= 6'h00;
      write_address_data_log_force[1842] <= 6'h00;
      write_address_data_log_force[1843] <= 6'h00;
      write_address_data_log_force[1844] <= 6'h00;
      write_address_data_log_force[1845] <= 6'h00;
      write_address_data_log_force[1846] <= 6'h00;
      write_address_data_log_force[1847] <= 6'h00;
      write_address_data_log_force[1848] <= 6'h00;
      write_address_data_log_force[1849] <= 6'h00;
      write_address_data_log_force[1850] <= 6'h00;
      write_address_data_log_force[1851] <= 6'h00;
      write_address_data_log_force[1852] <= 6'h00;
      write_address_data_log_force[1853] <= 6'h00;
      write_address_data_log_force[1854] <= 6'h00;
      write_address_data_log_force[1855] <= 6'h00;
      write_address_data_log_force[1856] <= 6'h00;
      write_address_data_log_force[1857] <= 6'h00;
      write_address_data_log_force[1858] <= 6'h00;
      write_address_data_log_force[1859] <= 6'h00;
      write_address_data_log_force[1860] <= 6'h00;
      write_address_data_log_force[1861] <= 6'h00;
      write_address_data_log_force[1862] <= 6'h00;
      write_address_data_log_force[1863] <= 6'h00;
      write_address_data_log_force[1864] <= 6'h00;
      write_address_data_log_force[1865] <= 6'h00;
      write_address_data_log_force[1866] <= 6'h00;
      write_address_data_log_force[1867] <= 6'h00;
      write_address_data_log_force[1868] <= 6'h00;
      write_address_data_log_force[1869] <= 6'h00;
      write_address_data_log_force[1870] <= 6'h00;
      write_address_data_log_force[1871] <= 6'h00;
      write_address_data_log_force[1872] <= 6'h00;
      write_address_data_log_force[1873] <= 6'h00;
      write_address_data_log_force[1874] <= 6'h00;
      write_address_data_log_force[1875] <= 6'h00;
      write_address_data_log_force[1876] <= 6'h00;
      write_address_data_log_force[1877] <= 6'h00;
      write_address_data_log_force[1878] <= 6'h00;
      write_address_data_log_force[1879] <= 6'h00;
      write_address_data_log_force[1880] <= 6'h00;
      write_address_data_log_force[1881] <= 6'h00;
      write_address_data_log_force[1882] <= 6'h00;
      write_address_data_log_force[1883] <= 6'h00;
      write_address_data_log_force[1884] <= 6'h00;
      write_address_data_log_force[1885] <= 6'h00;
      write_address_data_log_force[1886] <= 6'h00;
      write_address_data_log_force[1887] <= 6'h00;
      write_address_data_log_force[1888] <= 6'h00;
      write_address_data_log_force[1889] <= 6'h00;
      write_address_data_log_force[1890] <= 6'h00;
      write_address_data_log_force[1891] <= 6'h00;
      write_address_data_log_force[1892] <= 6'h00;
      write_address_data_log_force[1893] <= 6'h00;
      write_address_data_log_force[1894] <= 6'h00;
      write_address_data_log_force[1895] <= 6'h00;
      write_address_data_log_force[1896] <= 6'h00;
      write_address_data_log_force[1897] <= 6'h00;
      write_address_data_log_force[1898] <= 6'h00;
      write_address_data_log_force[1899] <= 6'h00;
      write_address_data_log_force[1900] <= 6'h00;
      write_address_data_log_force[1901] <= 6'h00;
      write_address_data_log_force[1902] <= 6'h00;
      write_address_data_log_force[1903] <= 6'h00;
      write_address_data_log_force[1904] <= 6'h00;
      write_address_data_log_force[1905] <= 6'h00;
      write_address_data_log_force[1906] <= 6'h00;
      write_address_data_log_force[1907] <= 6'h00;
      write_address_data_log_force[1908] <= 6'h00;
      write_address_data_log_force[1909] <= 6'h00;
      write_address_data_log_force[1910] <= 6'h00;
      write_address_data_log_force[1911] <= 6'h00;
      write_address_data_log_force[1912] <= 6'h00;
      write_address_data_log_force[1913] <= 6'h00;
      write_address_data_log_force[1914] <= 6'h00;
      write_address_data_log_force[1915] <= 6'h00;
      write_address_data_log_force[1916] <= 6'h00;
      write_address_data_log_force[1917] <= 6'h00;
      write_address_data_log_force[1918] <= 6'h00;
      write_address_data_log_force[1919] <= 6'h00;
      write_address_data_log_force[1920] <= 6'h00;
      write_address_data_log_force[1921] <= 6'h00;
      write_address_data_log_force[1922] <= 6'h00;
      write_address_data_log_force[1923] <= 6'h00;
      write_address_data_log_force[1924] <= 6'h00;
      write_address_data_log_force[1925] <= 6'h00;
      write_address_data_log_force[1926] <= 6'h00;
      write_address_data_log_force[1927] <= 6'h00;
      write_address_data_log_force[1928] <= 6'h00;
      write_address_data_log_force[1929] <= 6'h00;
      write_address_data_log_force[1930] <= 6'h00;
      write_address_data_log_force[1931] <= 6'h00;
      write_address_data_log_force[1932] <= 6'h00;
      write_address_data_log_force[1933] <= 6'h00;
      write_address_data_log_force[1934] <= 6'h00;
      write_address_data_log_force[1935] <= 6'h00;
      write_address_data_log_force[1936] <= 6'h00;
      write_address_data_log_force[1937] <= 6'h00;
      write_address_data_log_force[1938] <= 6'h00;
      write_address_data_log_force[1939] <= 6'h00;
      write_address_data_log_force[1940] <= 6'h00;
      write_address_data_log_force[1941] <= 6'h00;
      write_address_data_log_force[1942] <= 6'h00;
      write_address_data_log_force[1943] <= 6'h00;
      write_address_data_log_force[1944] <= 6'h00;
      write_address_data_log_force[1945] <= 6'h00;
      write_address_data_log_force[1946] <= 6'h00;
      write_address_data_log_force[1947] <= 6'h00;
      write_address_data_log_force[1948] <= 6'h00;
      write_address_data_log_force[1949] <= 6'h00;
      write_address_data_log_force[1950] <= 6'h00;
      write_address_data_log_force[1951] <= 6'h00;
      write_address_data_log_force[1952] <= 6'h00;
      write_address_data_log_force[1953] <= 6'h00;
      write_address_data_log_force[1954] <= 6'h00;
      write_address_data_log_force[1955] <= 6'h00;
      write_address_data_log_force[1956] <= 6'h00;
      write_address_data_log_force[1957] <= 6'h00;
      write_address_data_log_force[1958] <= 6'h00;
      write_address_data_log_force[1959] <= 6'h00;
      write_address_data_log_force[1960] <= 6'h00;
      write_address_data_log_force[1961] <= 6'h00;
      write_address_data_log_force[1962] <= 6'h00;
      write_address_data_log_force[1963] <= 6'h00;
      write_address_data_log_force[1964] <= 6'h00;
      write_address_data_log_force[1965] <= 6'h00;
      write_address_data_log_force[1966] <= 6'h00;
      write_address_data_log_force[1967] <= 6'h00;
      write_address_data_log_force[1968] <= 6'h00;
      write_address_data_log_force[1969] <= 6'h00;
      write_address_data_log_force[1970] <= 6'h00;
      write_address_data_log_force[1971] <= 6'h00;
      write_address_data_log_force[1972] <= 6'h00;
      write_address_data_log_force[1973] <= 6'h00;
      write_address_data_log_force[1974] <= 6'h00;
      write_address_data_log_force[1975] <= 6'h00;
      write_address_data_log_force[1976] <= 6'h00;
      write_address_data_log_force[1977] <= 6'h00;
      write_address_data_log_force[1978] <= 6'h00;
      write_address_data_log_force[1979] <= 6'h00;
      write_address_data_log_force[1980] <= 6'h00;
      write_address_data_log_force[1981] <= 6'h00;
      write_address_data_log_force[1982] <= 6'h00;
      write_address_data_log_force[1983] <= 6'h00;
      write_address_data_log_force[1984] <= 6'h00;
      write_address_data_log_force[1985] <= 6'h00;
      write_address_data_log_force[1986] <= 6'h00;
      write_address_data_log_force[1987] <= 6'h00;
      write_address_data_log_force[1988] <= 6'h00;
      write_address_data_log_force[1989] <= 6'h00;
      write_address_data_log_force[1990] <= 6'h00;
      write_address_data_log_force[1991] <= 6'h00;
      write_address_data_log_force[1992] <= 6'h00;
      write_address_data_log_force[1993] <= 6'h00;
      write_address_data_log_force[1994] <= 6'h00;
      write_address_data_log_force[1995] <= 6'h00;
      write_address_data_log_force[1996] <= 6'h00;
      write_address_data_log_force[1997] <= 6'h00;
      write_address_data_log_force[1998] <= 6'h00;
      write_address_data_log_force[1999] <= 6'h00;
      write_address_data_log_force[2000] <= 6'h00;
      write_address_data_log_force[2001] <= 6'h00;
      write_address_data_log_force[2002] <= 6'h00;
      write_address_data_log_force[2003] <= 6'h00;
      write_address_data_log_force[2004] <= 6'h00;
      write_address_data_log_force[2005] <= 6'h00;
      write_address_data_log_force[2006] <= 6'h00;
      write_address_data_log_force[2007] <= 6'h00;
      write_address_data_log_force[2008] <= 6'h00;
      write_address_data_log_force[2009] <= 6'h00;
      write_address_data_log_force[2010] <= 6'h00;
      write_address_data_log_force[2011] <= 6'h00;
      write_address_data_log_force[2012] <= 6'h00;
      write_address_data_log_force[2013] <= 6'h00;
      write_address_data_log_force[2014] <= 6'h00;
      write_address_data_log_force[2015] <= 6'h00;
      write_address_data_log_force[2016] <= 6'h00;
      write_address_data_log_force[2017] <= 6'h00;
      write_address_data_log_force[2018] <= 6'h00;
      write_address_data_log_force[2019] <= 6'h00;
      write_address_data_log_force[2020] <= 6'h00;
      write_address_data_log_force[2021] <= 6'h00;
      write_address_data_log_force[2022] <= 6'h00;
      write_address_data_log_force[2023] <= 6'h00;
      write_address_data_log_force[2024] <= 6'h00;
      write_address_data_log_force[2025] <= 6'h00;
      write_address_data_log_force[2026] <= 6'h00;
      write_address_data_log_force[2027] <= 6'h00;
      write_address_data_log_force[2028] <= 6'h00;
      write_address_data_log_force[2029] <= 6'h00;
      write_address_data_log_force[2030] <= 6'h00;
      write_address_data_log_force[2031] <= 6'h00;
      write_address_data_log_force[2032] <= 6'h00;
      write_address_data_log_force[2033] <= 6'h00;
      write_address_data_log_force[2034] <= 6'h00;
      write_address_data_log_force[2035] <= 6'h00;
      write_address_data_log_force[2036] <= 6'h00;
      write_address_data_log_force[2037] <= 6'h00;
      write_address_data_log_force[2038] <= 6'h00;
      write_address_data_log_force[2039] <= 6'h00;
      write_address_data_log_force[2040] <= 6'h00;
      write_address_data_log_force[2041] <= 6'h00;
      write_address_data_log_force[2042] <= 6'h00;
      write_address_data_log_force[2043] <= 6'h00;
      write_address_data_log_force[2044] <= 6'h00;
      write_address_data_log_force[2045] <= 6'h00;
      write_address_data_log_force[2046] <= 6'h00;
      write_address_data_log_force[2047] <= 6'h00;
      write_address_data_log_force[2048] <= 6'h00;
      write_address_data_log_force[2049] <= 6'h00;
      write_address_data_log_force[2050] <= 6'h00;
      write_address_data_log_force[2051] <= 6'h00;
      write_address_data_log_force[2052] <= 6'h00;
      write_address_data_log_force[2053] <= 6'h00;
      write_address_data_log_force[2054] <= 6'h00;
      write_address_data_log_force[2055] <= 6'h00;
      write_address_data_log_force[2056] <= 6'h00;
      write_address_data_log_force[2057] <= 6'h00;
      write_address_data_log_force[2058] <= 6'h00;
      write_address_data_log_force[2059] <= 6'h00;
      write_address_data_log_force[2060] <= 6'h00;
      write_address_data_log_force[2061] <= 6'h00;
      write_address_data_log_force[2062] <= 6'h00;
      write_address_data_log_force[2063] <= 6'h00;
      write_address_data_log_force[2064] <= 6'h00;
      write_address_data_log_force[2065] <= 6'h00;
      write_address_data_log_force[2066] <= 6'h00;
      write_address_data_log_force[2067] <= 6'h00;
      write_address_data_log_force[2068] <= 6'h00;
      write_address_data_log_force[2069] <= 6'h00;
      write_address_data_log_force[2070] <= 6'h00;
      write_address_data_log_force[2071] <= 6'h00;
      write_address_data_log_force[2072] <= 6'h00;
      write_address_data_log_force[2073] <= 6'h00;
      write_address_data_log_force[2074] <= 6'h00;
      write_address_data_log_force[2075] <= 6'h00;
      write_address_data_log_force[2076] <= 6'h00;
      write_address_data_log_force[2077] <= 6'h00;
      write_address_data_log_force[2078] <= 6'h00;
      write_address_data_log_force[2079] <= 6'h00;
      write_address_data_log_force[2080] <= 6'h00;
      write_address_data_log_force[2081] <= 6'h00;
      write_address_data_log_force[2082] <= 6'h00;
      write_address_data_log_force[2083] <= 6'h00;
      write_address_data_log_force[2084] <= 6'h00;
      write_address_data_log_force[2085] <= 6'h00;
      write_address_data_log_force[2086] <= 6'h00;
      write_address_data_log_force[2087] <= 6'h00;
      write_address_data_log_force[2088] <= 6'h00;
      write_address_data_log_force[2089] <= 6'h00;
      write_address_data_log_force[2090] <= 6'h00;
      write_address_data_log_force[2091] <= 6'h00;
      write_address_data_log_force[2092] <= 6'h00;
      write_address_data_log_force[2093] <= 6'h00;
      write_address_data_log_force[2094] <= 6'h00;
      write_address_data_log_force[2095] <= 6'h00;
      write_address_data_log_force[2096] <= 6'h00;
      write_address_data_log_force[2097] <= 6'h00;
      write_address_data_log_force[2098] <= 6'h00;
      write_address_data_log_force[2099] <= 6'h00;
      write_address_data_log_force[2100] <= 6'h00;
      write_address_data_log_force[2101] <= 6'h00;
      write_address_data_log_force[2102] <= 6'h00;
      write_address_data_log_force[2103] <= 6'h00;
      write_address_data_log_force[2104] <= 6'h00;
      write_address_data_log_force[2105] <= 6'h00;
      write_address_data_log_force[2106] <= 6'h00;
      write_address_data_log_force[2107] <= 6'h00;
      write_address_data_log_force[2108] <= 6'h00;
      write_address_data_log_force[2109] <= 6'h00;
      write_address_data_log_force[2110] <= 6'h00;
      write_address_data_log_force[2111] <= 6'h00;
      write_address_data_log_force[2112] <= 6'h00;
      write_address_data_log_force[2113] <= 6'h00;
      write_address_data_log_force[2114] <= 6'h00;
      write_address_data_log_force[2115] <= 6'h00;
      write_address_data_log_force[2116] <= 6'h00;
      write_address_data_log_force[2117] <= 6'h00;
      write_address_data_log_force[2118] <= 6'h00;
      write_address_data_log_force[2119] <= 6'h00;
      write_address_data_log_force[2120] <= 6'h00;
      write_address_data_log_force[2121] <= 6'h00;
      write_address_data_log_force[2122] <= 6'h00;
      write_address_data_log_force[2123] <= 6'h00;
      write_address_data_log_force[2124] <= 6'h00;
      write_address_data_log_force[2125] <= 6'h00;
      write_address_data_log_force[2126] <= 6'h00;
      write_address_data_log_force[2127] <= 6'h00;
      write_address_data_log_force[2128] <= 6'h00;
      write_address_data_log_force[2129] <= 6'h00;
      write_address_data_log_force[2130] <= 6'h00;
      write_address_data_log_force[2131] <= 6'h00;
      write_address_data_log_force[2132] <= 6'h00;
      write_address_data_log_force[2133] <= 6'h00;
      write_address_data_log_force[2134] <= 6'h00;
      write_address_data_log_force[2135] <= 6'h00;
      write_address_data_log_force[2136] <= 6'h00;
      write_address_data_log_force[2137] <= 6'h00;
      write_address_data_log_force[2138] <= 6'h00;
      write_address_data_log_force[2139] <= 6'h00;
      write_address_data_log_force[2140] <= 6'h00;
      write_address_data_log_force[2141] <= 6'h00;
      write_address_data_log_force[2142] <= 6'h00;
      write_address_data_log_force[2143] <= 6'h00;
      write_address_data_log_force[2144] <= 6'h00;
      write_address_data_log_force[2145] <= 6'h00;
      write_address_data_log_force[2146] <= 6'h00;
      write_address_data_log_force[2147] <= 6'h00;
      write_address_data_log_force[2148] <= 6'h00;
      write_address_data_log_force[2149] <= 6'h00;
      write_address_data_log_force[2150] <= 6'h00;
      write_address_data_log_force[2151] <= 6'h00;
      write_address_data_log_force[2152] <= 6'h00;
      write_address_data_log_force[2153] <= 6'h00;
      write_address_data_log_force[2154] <= 6'h00;
      write_address_data_log_force[2155] <= 6'h00;
      write_address_data_log_force[2156] <= 6'h00;
      write_address_data_log_force[2157] <= 6'h00;
      write_address_data_log_force[2158] <= 6'h00;
      write_address_data_log_force[2159] <= 6'h00;
      write_address_data_log_force[2160] <= 6'h00;
      write_address_data_log_force[2161] <= 6'h00;
      write_address_data_log_force[2162] <= 6'h00;
      write_address_data_log_force[2163] <= 6'h00;
      write_address_data_log_force[2164] <= 6'h00;
      write_address_data_log_force[2165] <= 6'h00;
      write_address_data_log_force[2166] <= 6'h00;
      write_address_data_log_force[2167] <= 6'h00;
      write_address_data_log_force[2168] <= 6'h00;
      write_address_data_log_force[2169] <= 6'h00;
      write_address_data_log_force[2170] <= 6'h00;
      write_address_data_log_force[2171] <= 6'h00;
      write_address_data_log_force[2172] <= 6'h00;
      write_address_data_log_force[2173] <= 6'h00;
      write_address_data_log_force[2174] <= 6'h00;
      write_address_data_log_force[2175] <= 6'h00;
      write_address_data_log_force[2176] <= 6'h00;
      write_address_data_log_force[2177] <= 6'h00;
      write_address_data_log_force[2178] <= 6'h00;
      write_address_data_log_force[2179] <= 6'h00;
      write_address_data_log_force[2180] <= 6'h00;
      write_address_data_log_force[2181] <= 6'h00;
      write_address_data_log_force[2182] <= 6'h00;
      write_address_data_log_force[2183] <= 6'h00;
      write_address_data_log_force[2184] <= 6'h00;
      write_address_data_log_force[2185] <= 6'h00;
      write_address_data_log_force[2186] <= 6'h00;
      write_address_data_log_force[2187] <= 6'h00;
      write_address_data_log_force[2188] <= 6'h00;
      write_address_data_log_force[2189] <= 6'h00;
      write_address_data_log_force[2190] <= 6'h00;
      write_address_data_log_force[2191] <= 6'h00;
      write_address_data_log_force[2192] <= 6'h00;
      write_address_data_log_force[2193] <= 6'h00;
      write_address_data_log_force[2194] <= 6'h00;
      write_address_data_log_force[2195] <= 6'h00;
      write_address_data_log_force[2196] <= 6'h00;
      write_address_data_log_force[2197] <= 6'h00;
      write_address_data_log_force[2198] <= 6'h00;
      write_address_data_log_force[2199] <= 6'h00;
      write_address_data_log_force[2200] <= 6'h00;
      write_address_data_log_force[2201] <= 6'h00;
      write_address_data_log_force[2202] <= 6'h00;
      write_address_data_log_force[2203] <= 6'h00;
      write_address_data_log_force[2204] <= 6'h00;
      write_address_data_log_force[2205] <= 6'h00;
      write_address_data_log_force[2206] <= 6'h00;
      write_address_data_log_force[2207] <= 6'h00;
      write_address_data_log_force[2208] <= 6'h00;
      write_address_data_log_force[2209] <= 6'h00;
      write_address_data_log_force[2210] <= 6'h00;
      write_address_data_log_force[2211] <= 6'h00;
      write_address_data_log_force[2212] <= 6'h00;
      write_address_data_log_force[2213] <= 6'h00;
      write_address_data_log_force[2214] <= 6'h00;
      write_address_data_log_force[2215] <= 6'h00;
      write_address_data_log_force[2216] <= 6'h00;
      write_address_data_log_force[2217] <= 6'h00;
      write_address_data_log_force[2218] <= 6'h00;
      write_address_data_log_force[2219] <= 6'h00;
      write_address_data_log_force[2220] <= 6'h00;
      write_address_data_log_force[2221] <= 6'h00;
      write_address_data_log_force[2222] <= 6'h00;
      write_address_data_log_force[2223] <= 6'h00;
      write_address_data_log_force[2224] <= 6'h00;
      write_address_data_log_force[2225] <= 6'h00;
      write_address_data_log_force[2226] <= 6'h00;
      write_address_data_log_force[2227] <= 6'h00;
      write_address_data_log_force[2228] <= 6'h00;
      write_address_data_log_force[2229] <= 6'h00;
      write_address_data_log_force[2230] <= 6'h00;
      write_address_data_log_force[2231] <= 6'h00;
      write_address_data_log_force[2232] <= 6'h00;
      write_address_data_log_force[2233] <= 6'h00;
      write_address_data_log_force[2234] <= 6'h00;
      write_address_data_log_force[2235] <= 6'h00;
      write_address_data_log_force[2236] <= 6'h00;
      write_address_data_log_force[2237] <= 6'h00;
      write_address_data_log_force[2238] <= 6'h00;
      write_address_data_log_force[2239] <= 6'h00;
      write_address_data_log_force[2240] <= 6'h00;
      write_address_data_log_force[2241] <= 6'h00;
      write_address_data_log_force[2242] <= 6'h00;
      write_address_data_log_force[2243] <= 6'h00;
      write_address_data_log_force[2244] <= 6'h00;
      write_address_data_log_force[2245] <= 6'h00;
      write_address_data_log_force[2246] <= 6'h00;
      write_address_data_log_force[2247] <= 6'h00;
      write_address_data_log_force[2248] <= 6'h00;
      write_address_data_log_force[2249] <= 6'h00;
      write_address_data_log_force[2250] <= 6'h00;
      write_address_data_log_force[2251] <= 6'h00;
      write_address_data_log_force[2252] <= 6'h00;
      write_address_data_log_force[2253] <= 6'h00;
      write_address_data_log_force[2254] <= 6'h00;
      write_address_data_log_force[2255] <= 6'h00;
      write_address_data_log_force[2256] <= 6'h00;
      write_address_data_log_force[2257] <= 6'h00;
      write_address_data_log_force[2258] <= 6'h00;
      write_address_data_log_force[2259] <= 6'h00;
      write_address_data_log_force[2260] <= 6'h00;
      write_address_data_log_force[2261] <= 6'h00;
      write_address_data_log_force[2262] <= 6'h00;
      write_address_data_log_force[2263] <= 6'h00;
      write_address_data_log_force[2264] <= 6'h00;
      write_address_data_log_force[2265] <= 6'h00;
      write_address_data_log_force[2266] <= 6'h00;
      write_address_data_log_force[2267] <= 6'h00;
      write_address_data_log_force[2268] <= 6'h00;
      write_address_data_log_force[2269] <= 6'h00;
      write_address_data_log_force[2270] <= 6'h00;
      write_address_data_log_force[2271] <= 6'h00;
      write_address_data_log_force[2272] <= 6'h00;
      write_address_data_log_force[2273] <= 6'h00;
      write_address_data_log_force[2274] <= 6'h00;
      write_address_data_log_force[2275] <= 6'h00;
      write_address_data_log_force[2276] <= 6'h00;
      write_address_data_log_force[2277] <= 6'h00;
      write_address_data_log_force[2278] <= 6'h00;
      write_address_data_log_force[2279] <= 6'h00;
      write_address_data_log_force[2280] <= 6'h00;
      write_address_data_log_force[2281] <= 6'h00;
      write_address_data_log_force[2282] <= 6'h00;
      write_address_data_log_force[2283] <= 6'h00;
      write_address_data_log_force[2284] <= 6'h00;
      write_address_data_log_force[2285] <= 6'h00;
      write_address_data_log_force[2286] <= 6'h00;
      write_address_data_log_force[2287] <= 6'h00;
      write_address_data_log_force[2288] <= 6'h00;
      write_address_data_log_force[2289] <= 6'h00;
      write_address_data_log_force[2290] <= 6'h00;
      write_address_data_log_force[2291] <= 6'h00;
      write_address_data_log_force[2292] <= 6'h00;
      write_address_data_log_force[2293] <= 6'h00;
      write_address_data_log_force[2294] <= 6'h00;
      write_address_data_log_force[2295] <= 6'h00;
      write_address_data_log_force[2296] <= 6'h00;
      write_address_data_log_force[2297] <= 6'h00;
      write_address_data_log_force[2298] <= 6'h00;
      write_address_data_log_force[2299] <= 6'h00;
      write_address_data_log_force[2300] <= 6'h00;
      write_address_data_log_force[2301] <= 6'h00;
      write_address_data_log_force[2302] <= 6'h00;
      write_address_data_log_force[2303] <= 6'h00;
      write_address_data_log_force[2304] <= 6'h00;
      write_address_data_log_force[2305] <= 6'h00;
      write_address_data_log_force[2306] <= 6'h00;
      write_address_data_log_force[2307] <= 6'h00;
      write_address_data_log_force[2308] <= 6'h00;
      write_address_data_log_force[2309] <= 6'h00;
      write_address_data_log_force[2310] <= 6'h00;
      write_address_data_log_force[2311] <= 6'h00;
      write_address_data_log_force[2312] <= 6'h00;
      write_address_data_log_force[2313] <= 6'h00;
      write_address_data_log_force[2314] <= 6'h00;
      write_address_data_log_force[2315] <= 6'h00;
      write_address_data_log_force[2316] <= 6'h00;
      write_address_data_log_force[2317] <= 6'h00;
      write_address_data_log_force[2318] <= 6'h00;
      write_address_data_log_force[2319] <= 6'h00;
      write_address_data_log_force[2320] <= 6'h00;
      write_address_data_log_force[2321] <= 6'h00;
      write_address_data_log_force[2322] <= 6'h00;
      write_address_data_log_force[2323] <= 6'h00;
      write_address_data_log_force[2324] <= 6'h00;
      write_address_data_log_force[2325] <= 6'h00;
      write_address_data_log_force[2326] <= 6'h00;
      write_address_data_log_force[2327] <= 6'h00;
      write_address_data_log_force[2328] <= 6'h00;
      write_address_data_log_force[2329] <= 6'h00;
      write_address_data_log_force[2330] <= 6'h00;
      write_address_data_log_force[2331] <= 6'h00;
      write_address_data_log_force[2332] <= 6'h00;
      write_address_data_log_force[2333] <= 6'h00;
      write_address_data_log_force[2334] <= 6'h00;
      write_address_data_log_force[2335] <= 6'h00;
      write_address_data_log_force[2336] <= 6'h00;
      write_address_data_log_force[2337] <= 6'h00;
      write_address_data_log_force[2338] <= 6'h00;
      write_address_data_log_force[2339] <= 6'h00;
      write_address_data_log_force[2340] <= 6'h00;
      write_address_data_log_force[2341] <= 6'h00;
      write_address_data_log_force[2342] <= 6'h00;
      write_address_data_log_force[2343] <= 6'h00;
      write_address_data_log_force[2344] <= 6'h00;
      write_address_data_log_force[2345] <= 6'h00;
      write_address_data_log_force[2346] <= 6'h00;
      write_address_data_log_force[2347] <= 6'h00;
      write_address_data_log_force[2348] <= 6'h00;
      write_address_data_log_force[2349] <= 6'h00;
      write_address_data_log_force[2350] <= 6'h00;
      write_address_data_log_force[2351] <= 6'h00;
      write_address_data_log_force[2352] <= 6'h00;
      write_address_data_log_force[2353] <= 6'h00;
      write_address_data_log_force[2354] <= 6'h00;
      write_address_data_log_force[2355] <= 6'h00;
      write_address_data_log_force[2356] <= 6'h00;
      write_address_data_log_force[2357] <= 6'h00;
      write_address_data_log_force[2358] <= 6'h00;
      write_address_data_log_force[2359] <= 6'h00;
      write_address_data_log_force[2360] <= 6'h00;
      write_address_data_log_force[2361] <= 6'h00;
      write_address_data_log_force[2362] <= 6'h00;
      write_address_data_log_force[2363] <= 6'h00;
      write_address_data_log_force[2364] <= 6'h00;
      write_address_data_log_force[2365] <= 6'h00;
      write_address_data_log_force[2366] <= 6'h00;
      write_address_data_log_force[2367] <= 6'h00;
      write_address_data_log_force[2368] <= 6'h00;
      write_address_data_log_force[2369] <= 6'h00;
      write_address_data_log_force[2370] <= 6'h00;
      write_address_data_log_force[2371] <= 6'h00;
      write_address_data_log_force[2372] <= 6'h00;
      write_address_data_log_force[2373] <= 6'h00;
      write_address_data_log_force[2374] <= 6'h00;
      write_address_data_log_force[2375] <= 6'h00;
      write_address_data_log_force[2376] <= 6'h00;
      write_address_data_log_force[2377] <= 6'h00;
      write_address_data_log_force[2378] <= 6'h00;
      write_address_data_log_force[2379] <= 6'h00;
      write_address_data_log_force[2380] <= 6'h00;
      write_address_data_log_force[2381] <= 6'h00;
      write_address_data_log_force[2382] <= 6'h00;
      write_address_data_log_force[2383] <= 6'h00;
      write_address_data_log_force[2384] <= 6'h00;
      write_address_data_log_force[2385] <= 6'h00;
      write_address_data_log_force[2386] <= 6'h00;
      write_address_data_log_force[2387] <= 6'h00;
      write_address_data_log_force[2388] <= 6'h00;
      write_address_data_log_force[2389] <= 6'h00;
      write_address_data_log_force[2390] <= 6'h00;
      write_address_data_log_force[2391] <= 6'h00;
      write_address_data_log_force[2392] <= 6'h00;
      write_address_data_log_force[2393] <= 6'h00;
      write_address_data_log_force[2394] <= 6'h00;
      write_address_data_log_force[2395] <= 6'h00;
      write_address_data_log_force[2396] <= 6'h00;
      write_address_data_log_force[2397] <= 6'h00;
      write_address_data_log_force[2398] <= 6'h00;
      write_address_data_log_force[2399] <= 6'h00;
      write_address_data_log_force[2400] <= 6'h00;
      write_address_data_log_force[2401] <= 6'h00;
      write_address_data_log_force[2402] <= 6'h00;
      write_address_data_log_force[2403] <= 6'h00;
      write_address_data_log_force[2404] <= 6'h00;
      write_address_data_log_force[2405] <= 6'h00;
      write_address_data_log_force[2406] <= 6'h00;
      write_address_data_log_force[2407] <= 6'h00;
      write_address_data_log_force[2408] <= 6'h00;
      write_address_data_log_force[2409] <= 6'h00;
      write_address_data_log_force[2410] <= 6'h00;
      write_address_data_log_force[2411] <= 6'h00;
      write_address_data_log_force[2412] <= 6'h00;
      write_address_data_log_force[2413] <= 6'h00;
      write_address_data_log_force[2414] <= 6'h00;
      write_address_data_log_force[2415] <= 6'h00;
      write_address_data_log_force[2416] <= 6'h00;
      write_address_data_log_force[2417] <= 6'h00;
      write_address_data_log_force[2418] <= 6'h00;
      write_address_data_log_force[2419] <= 6'h00;
      write_address_data_log_force[2420] <= 6'h00;
      write_address_data_log_force[2421] <= 6'h00;
      write_address_data_log_force[2422] <= 6'h00;
      write_address_data_log_force[2423] <= 6'h00;
      write_address_data_log_force[2424] <= 6'h00;
      write_address_data_log_force[2425] <= 6'h00;
      write_address_data_log_force[2426] <= 6'h00;
      write_address_data_log_force[2427] <= 6'h00;
      write_address_data_log_force[2428] <= 6'h00;
      write_address_data_log_force[2429] <= 6'h00;
      write_address_data_log_force[2430] <= 6'h00;
      write_address_data_log_force[2431] <= 6'h00;
      write_address_data_log_force[2432] <= 6'h00;
      write_address_data_log_force[2433] <= 6'h00;
      write_address_data_log_force[2434] <= 6'h00;
      write_address_data_log_force[2435] <= 6'h00;
      write_address_data_log_force[2436] <= 6'h00;
      write_address_data_log_force[2437] <= 6'h00;
      write_address_data_log_force[2438] <= 6'h00;
      write_address_data_log_force[2439] <= 6'h00;
      write_address_data_log_force[2440] <= 6'h00;
      write_address_data_log_force[2441] <= 6'h00;
      write_address_data_log_force[2442] <= 6'h00;
      write_address_data_log_force[2443] <= 6'h00;
      write_address_data_log_force[2444] <= 6'h00;
      write_address_data_log_force[2445] <= 6'h00;
      write_address_data_log_force[2446] <= 6'h00;
      write_address_data_log_force[2447] <= 6'h00;
      write_address_data_log_force[2448] <= 6'h00;
      write_address_data_log_force[2449] <= 6'h00;
      write_address_data_log_force[2450] <= 6'h00;
      write_address_data_log_force[2451] <= 6'h00;
      write_address_data_log_force[2452] <= 6'h00;
      write_address_data_log_force[2453] <= 6'h00;
      write_address_data_log_force[2454] <= 6'h00;
      write_address_data_log_force[2455] <= 6'h00;
      write_address_data_log_force[2456] <= 6'h00;
      write_address_data_log_force[2457] <= 6'h00;
      write_address_data_log_force[2458] <= 6'h00;
      write_address_data_log_force[2459] <= 6'h00;
      write_address_data_log_force[2460] <= 6'h00;
      write_address_data_log_force[2461] <= 6'h00;
      write_address_data_log_force[2462] <= 6'h00;
      write_address_data_log_force[2463] <= 6'h00;
      write_address_data_log_force[2464] <= 6'h00;
      write_address_data_log_force[2465] <= 6'h00;
      write_address_data_log_force[2466] <= 6'h00;
      write_address_data_log_force[2467] <= 6'h00;
      write_address_data_log_force[2468] <= 6'h00;
      write_address_data_log_force[2469] <= 6'h00;
      write_address_data_log_force[2470] <= 6'h00;
      write_address_data_log_force[2471] <= 6'h00;
      write_address_data_log_force[2472] <= 6'h00;
      write_address_data_log_force[2473] <= 6'h00;
      write_address_data_log_force[2474] <= 6'h00;
      write_address_data_log_force[2475] <= 6'h00;
      write_address_data_log_force[2476] <= 6'h00;
      write_address_data_log_force[2477] <= 6'h00;
      write_address_data_log_force[2478] <= 6'h00;
      write_address_data_log_force[2479] <= 6'h00;
      write_address_data_log_force[2480] <= 6'h00;
      write_address_data_log_force[2481] <= 6'h00;
      write_address_data_log_force[2482] <= 6'h00;
      write_address_data_log_force[2483] <= 6'h00;
      write_address_data_log_force[2484] <= 6'h00;
      write_address_data_log_force[2485] <= 6'h00;
      write_address_data_log_force[2486] <= 6'h00;
      write_address_data_log_force[2487] <= 6'h00;
      write_address_data_log_force[2488] <= 6'h00;
      write_address_data_log_force[2489] <= 6'h00;
      write_address_data_log_force[2490] <= 6'h00;
      write_address_data_log_force[2491] <= 6'h00;
      write_address_data_log_force[2492] <= 6'h00;
      write_address_data_log_force[2493] <= 6'h00;
      write_address_data_log_force[2494] <= 6'h00;
      write_address_data_log_force[2495] <= 6'h00;
      write_address_data_log_force[2496] <= 6'h00;
      write_address_data_log_force[2497] <= 6'h00;
      write_address_data_log_force[2498] <= 6'h00;
      write_address_data_log_force[2499] <= 6'h00;
      write_address_data_log_force[2500] <= 6'h00;
      write_address_data_log_force[2501] <= 6'h00;
      write_address_data_log_force[2502] <= 6'h00;
      write_address_data_log_force[2503] <= 6'h00;
      write_address_data_log_force[2504] <= 6'h00;
      write_address_data_log_force[2505] <= 6'h00;
      write_address_data_log_force[2506] <= 6'h00;
      write_address_data_log_force[2507] <= 6'h00;
      write_address_data_log_force[2508] <= 6'h00;
      write_address_data_log_force[2509] <= 6'h00;
      write_address_data_log_force[2510] <= 6'h00;
      write_address_data_log_force[2511] <= 6'h00;
      write_address_data_log_force[2512] <= 6'h00;
      write_address_data_log_force[2513] <= 6'h00;
      write_address_data_log_force[2514] <= 6'h00;
      write_address_data_log_force[2515] <= 6'h00;
      write_address_data_log_force[2516] <= 6'h00;
      write_address_data_log_force[2517] <= 6'h00;
      write_address_data_log_force[2518] <= 6'h00;
      write_address_data_log_force[2519] <= 6'h00;
      write_address_data_log_force[2520] <= 6'h00;
      write_address_data_log_force[2521] <= 6'h00;
      write_address_data_log_force[2522] <= 6'h00;
      write_address_data_log_force[2523] <= 6'h00;
      write_address_data_log_force[2524] <= 6'h00;
      write_address_data_log_force[2525] <= 6'h00;
      write_address_data_log_force[2526] <= 6'h00;
      write_address_data_log_force[2527] <= 6'h00;
      write_address_data_log_force[2528] <= 6'h00;
      write_address_data_log_force[2529] <= 6'h00;
      write_address_data_log_force[2530] <= 6'h00;
      write_address_data_log_force[2531] <= 6'h00;
      write_address_data_log_force[2532] <= 6'h00;
      write_address_data_log_force[2533] <= 6'h00;
      write_address_data_log_force[2534] <= 6'h00;
      write_address_data_log_force[2535] <= 6'h00;
      write_address_data_log_force[2536] <= 6'h00;
      write_address_data_log_force[2537] <= 6'h00;
      write_address_data_log_force[2538] <= 6'h00;
      write_address_data_log_force[2539] <= 6'h00;
      write_address_data_log_force[2540] <= 6'h00;
      write_address_data_log_force[2541] <= 6'h00;
      write_address_data_log_force[2542] <= 6'h00;
      write_address_data_log_force[2543] <= 6'h00;
      write_address_data_log_force[2544] <= 6'h00;
      write_address_data_log_force[2545] <= 6'h00;
      write_address_data_log_force[2546] <= 6'h00;
      write_address_data_log_force[2547] <= 6'h00;
      write_address_data_log_force[2548] <= 6'h00;
      write_address_data_log_force[2549] <= 6'h00;
      write_address_data_log_force[2550] <= 6'h00;
      write_address_data_log_force[2551] <= 6'h00;
      write_address_data_log_force[2552] <= 6'h00;
      write_address_data_log_force[2553] <= 6'h00;
      write_address_data_log_force[2554] <= 6'h00;
      write_address_data_log_force[2555] <= 6'h00;
      write_address_data_log_force[2556] <= 6'h00;
      write_address_data_log_force[2557] <= 6'h00;
      write_address_data_log_force[2558] <= 6'h00;
      write_address_data_log_force[2559] <= 6'h00;
      write_address_data_log_force[2560] <= 6'h00;
      write_address_data_log_force[2561] <= 6'h00;
      write_address_data_log_force[2562] <= 6'h00;
      write_address_data_log_force[2563] <= 6'h00;
      write_address_data_log_force[2564] <= 6'h00;
      write_address_data_log_force[2565] <= 6'h00;
      write_address_data_log_force[2566] <= 6'h00;
      write_address_data_log_force[2567] <= 6'h00;
      write_address_data_log_force[2568] <= 6'h00;
      write_address_data_log_force[2569] <= 6'h00;
      write_address_data_log_force[2570] <= 6'h00;
      write_address_data_log_force[2571] <= 6'h00;
      write_address_data_log_force[2572] <= 6'h00;
      write_address_data_log_force[2573] <= 6'h00;
      write_address_data_log_force[2574] <= 6'h00;
      write_address_data_log_force[2575] <= 6'h00;
      write_address_data_log_force[2576] <= 6'h00;
      write_address_data_log_force[2577] <= 6'h00;
      write_address_data_log_force[2578] <= 6'h00;
      write_address_data_log_force[2579] <= 6'h00;
      write_address_data_log_force[2580] <= 6'h00;
      write_address_data_log_force[2581] <= 6'h00;
      write_address_data_log_force[2582] <= 6'h00;
      write_address_data_log_force[2583] <= 6'h00;
      write_address_data_log_force[2584] <= 6'h00;
      write_address_data_log_force[2585] <= 6'h00;
      write_address_data_log_force[2586] <= 6'h00;
      write_address_data_log_force[2587] <= 6'h00;
      write_address_data_log_force[2588] <= 6'h00;
      write_address_data_log_force[2589] <= 6'h00;
      write_address_data_log_force[2590] <= 6'h00;
      write_address_data_log_force[2591] <= 6'h00;
      write_address_data_log_force[2592] <= 6'h00;
      write_address_data_log_force[2593] <= 6'h00;
      write_address_data_log_force[2594] <= 6'h00;
      write_address_data_log_force[2595] <= 6'h00;
      write_address_data_log_force[2596] <= 6'h00;
      write_address_data_log_force[2597] <= 6'h00;
      write_address_data_log_force[2598] <= 6'h00;
      write_address_data_log_force[2599] <= 6'h00;
      write_address_data_log_force[2600] <= 6'h00;
      write_address_data_log_force[2601] <= 6'h00;
      write_address_data_log_force[2602] <= 6'h00;
      write_address_data_log_force[2603] <= 6'h00;
      write_address_data_log_force[2604] <= 6'h00;
      write_address_data_log_force[2605] <= 6'h00;
      write_address_data_log_force[2606] <= 6'h00;
      write_address_data_log_force[2607] <= 6'h00;
      write_address_data_log_force[2608] <= 6'h00;
      write_address_data_log_force[2609] <= 6'h00;
      write_address_data_log_force[2610] <= 6'h00;
      write_address_data_log_force[2611] <= 6'h00;
      write_address_data_log_force[2612] <= 6'h00;
      write_address_data_log_force[2613] <= 6'h00;
      write_address_data_log_force[2614] <= 6'h00;
      write_address_data_log_force[2615] <= 6'h00;
      write_address_data_log_force[2616] <= 6'h00;
      write_address_data_log_force[2617] <= 6'h00;
      write_address_data_log_force[2618] <= 6'h00;
      write_address_data_log_force[2619] <= 6'h00;
      write_address_data_log_force[2620] <= 6'h00;
      write_address_data_log_force[2621] <= 6'h00;
      write_address_data_log_force[2622] <= 6'h00;
      write_address_data_log_force[2623] <= 6'h00;
      write_address_data_log_force[2624] <= 6'h00;
      write_address_data_log_force[2625] <= 6'h00;
      write_address_data_log_force[2626] <= 6'h00;
      write_address_data_log_force[2627] <= 6'h00;
      write_address_data_log_force[2628] <= 6'h00;
      write_address_data_log_force[2629] <= 6'h00;
      write_address_data_log_force[2630] <= 6'h00;
      write_address_data_log_force[2631] <= 6'h00;
      write_address_data_log_force[2632] <= 6'h00;
      write_address_data_log_force[2633] <= 6'h00;
      write_address_data_log_force[2634] <= 6'h00;
      write_address_data_log_force[2635] <= 6'h00;
      write_address_data_log_force[2636] <= 6'h00;
      write_address_data_log_force[2637] <= 6'h00;
      write_address_data_log_force[2638] <= 6'h00;
      write_address_data_log_force[2639] <= 6'h00;
      write_address_data_log_force[2640] <= 6'h00;
      write_address_data_log_force[2641] <= 6'h00;
      write_address_data_log_force[2642] <= 6'h00;
      write_address_data_log_force[2643] <= 6'h00;
      write_address_data_log_force[2644] <= 6'h00;
      write_address_data_log_force[2645] <= 6'h00;
      write_address_data_log_force[2646] <= 6'h00;
      write_address_data_log_force[2647] <= 6'h00;
      write_address_data_log_force[2648] <= 6'h00;
      write_address_data_log_force[2649] <= 6'h00;
      write_address_data_log_force[2650] <= 6'h00;
      write_address_data_log_force[2651] <= 6'h00;
      write_address_data_log_force[2652] <= 6'h00;
      write_address_data_log_force[2653] <= 6'h00;
      write_address_data_log_force[2654] <= 6'h00;
      write_address_data_log_force[2655] <= 6'h00;
      write_address_data_log_force[2656] <= 6'h00;
      write_address_data_log_force[2657] <= 6'h00;
      write_address_data_log_force[2658] <= 6'h00;
      write_address_data_log_force[2659] <= 6'h00;
      write_address_data_log_force[2660] <= 6'h00;
      write_address_data_log_force[2661] <= 6'h00;
      write_address_data_log_force[2662] <= 6'h00;
      write_address_data_log_force[2663] <= 6'h00;
      write_address_data_log_force[2664] <= 6'h00;
      write_address_data_log_force[2665] <= 6'h00;
      write_address_data_log_force[2666] <= 6'h00;
      write_address_data_log_force[2667] <= 6'h00;
      write_address_data_log_force[2668] <= 6'h00;
      write_address_data_log_force[2669] <= 6'h00;
      write_address_data_log_force[2670] <= 6'h00;
      write_address_data_log_force[2671] <= 6'h00;
      write_address_data_log_force[2672] <= 6'h00;
      write_address_data_log_force[2673] <= 6'h00;
      write_address_data_log_force[2674] <= 6'h00;
      write_address_data_log_force[2675] <= 6'h00;
      write_address_data_log_force[2676] <= 6'h00;
      write_address_data_log_force[2677] <= 6'h00;
      write_address_data_log_force[2678] <= 6'h00;
      write_address_data_log_force[2679] <= 6'h00;
      write_address_data_log_force[2680] <= 6'h00;
      write_address_data_log_force[2681] <= 6'h00;
      write_address_data_log_force[2682] <= 6'h00;
      write_address_data_log_force[2683] <= 6'h00;
      write_address_data_log_force[2684] <= 6'h00;
      write_address_data_log_force[2685] <= 6'h00;
      write_address_data_log_force[2686] <= 6'h00;
      write_address_data_log_force[2687] <= 6'h00;
      write_address_data_log_force[2688] <= 6'h00;
      write_address_data_log_force[2689] <= 6'h00;
      write_address_data_log_force[2690] <= 6'h00;
      write_address_data_log_force[2691] <= 6'h00;
      write_address_data_log_force[2692] <= 6'h00;
      write_address_data_log_force[2693] <= 6'h00;
      write_address_data_log_force[2694] <= 6'h00;
      write_address_data_log_force[2695] <= 6'h00;
      write_address_data_log_force[2696] <= 6'h00;
      write_address_data_log_force[2697] <= 6'h00;
      write_address_data_log_force[2698] <= 6'h00;
      write_address_data_log_force[2699] <= 6'h00;
      write_address_data_log_force[2700] <= 6'h00;
      write_address_data_log_force[2701] <= 6'h00;
      write_address_data_log_force[2702] <= 6'h00;
      write_address_data_log_force[2703] <= 6'h00;
      write_address_data_log_force[2704] <= 6'h00;
      write_address_data_log_force[2705] <= 6'h00;
      write_address_data_log_force[2706] <= 6'h00;
      write_address_data_log_force[2707] <= 6'h00;
      write_address_data_log_force[2708] <= 6'h00;
      write_address_data_log_force[2709] <= 6'h00;
      write_address_data_log_force[2710] <= 6'h00;
      write_address_data_log_force[2711] <= 6'h00;
      write_address_data_log_force[2712] <= 6'h00;
      write_address_data_log_force[2713] <= 6'h00;
      write_address_data_log_force[2714] <= 6'h00;
      write_address_data_log_force[2715] <= 6'h00;
      write_address_data_log_force[2716] <= 6'h00;
      write_address_data_log_force[2717] <= 6'h00;
      write_address_data_log_force[2718] <= 6'h00;
      write_address_data_log_force[2719] <= 6'h00;
      write_address_data_log_force[2720] <= 6'h00;
      write_address_data_log_force[2721] <= 6'h00;
      write_address_data_log_force[2722] <= 6'h00;
      write_address_data_log_force[2723] <= 6'h00;
      write_address_data_log_force[2724] <= 6'h00;
      write_address_data_log_force[2725] <= 6'h00;
      write_address_data_log_force[2726] <= 6'h00;
      write_address_data_log_force[2727] <= 6'h00;
      write_address_data_log_force[2728] <= 6'h00;
      write_address_data_log_force[2729] <= 6'h00;
      write_address_data_log_force[2730] <= 6'h00;
      write_address_data_log_force[2731] <= 6'h00;
      write_address_data_log_force[2732] <= 6'h00;
      write_address_data_log_force[2733] <= 6'h00;
      write_address_data_log_force[2734] <= 6'h00;
      write_address_data_log_force[2735] <= 6'h00;
      write_address_data_log_force[2736] <= 6'h00;
      write_address_data_log_force[2737] <= 6'h00;
      write_address_data_log_force[2738] <= 6'h00;
      write_address_data_log_force[2739] <= 6'h00;
      write_address_data_log_force[2740] <= 6'h00;
      write_address_data_log_force[2741] <= 6'h00;
      write_address_data_log_force[2742] <= 6'h00;
      write_address_data_log_force[2743] <= 6'h00;
      write_address_data_log_force[2744] <= 6'h00;
      write_address_data_log_force[2745] <= 6'h00;
      write_address_data_log_force[2746] <= 6'h00;
      write_address_data_log_force[2747] <= 6'h00;
      write_address_data_log_force[2748] <= 6'h00;
      write_address_data_log_force[2749] <= 6'h00;
      write_address_data_log_force[2750] <= 6'h00;
      write_address_data_log_force[2751] <= 6'h00;
      write_address_data_log_force[2752] <= 6'h00;
      write_address_data_log_force[2753] <= 6'h00;
      write_address_data_log_force[2754] <= 6'h00;
      write_address_data_log_force[2755] <= 6'h00;
      write_address_data_log_force[2756] <= 6'h00;
      write_address_data_log_force[2757] <= 6'h00;
      write_address_data_log_force[2758] <= 6'h00;
      write_address_data_log_force[2759] <= 6'h00;
      write_address_data_log_force[2760] <= 6'h00;
      write_address_data_log_force[2761] <= 6'h00;
      write_address_data_log_force[2762] <= 6'h00;
      write_address_data_log_force[2763] <= 6'h00;
      write_address_data_log_force[2764] <= 6'h00;
      write_address_data_log_force[2765] <= 6'h00;
      write_address_data_log_force[2766] <= 6'h00;
      write_address_data_log_force[2767] <= 6'h00;
      write_address_data_log_force[2768] <= 6'h00;
      write_address_data_log_force[2769] <= 6'h00;
      write_address_data_log_force[2770] <= 6'h00;
      write_address_data_log_force[2771] <= 6'h00;
      write_address_data_log_force[2772] <= 6'h00;
      write_address_data_log_force[2773] <= 6'h00;
      write_address_data_log_force[2774] <= 6'h00;
      write_address_data_log_force[2775] <= 6'h00;
      write_address_data_log_force[2776] <= 6'h00;
      write_address_data_log_force[2777] <= 6'h00;
      write_address_data_log_force[2778] <= 6'h00;
      write_address_data_log_force[2779] <= 6'h00;
      write_address_data_log_force[2780] <= 6'h00;
      write_address_data_log_force[2781] <= 6'h00;
      write_address_data_log_force[2782] <= 6'h00;
      write_address_data_log_force[2783] <= 6'h00;
      write_address_data_log_force[2784] <= 6'h00;
      write_address_data_log_force[2785] <= 6'h00;
      write_address_data_log_force[2786] <= 6'h00;
      write_address_data_log_force[2787] <= 6'h00;
      write_address_data_log_force[2788] <= 6'h00;
      write_address_data_log_force[2789] <= 6'h00;
      write_address_data_log_force[2790] <= 6'h00;
      write_address_data_log_force[2791] <= 6'h00;
      write_address_data_log_force[2792] <= 6'h00;
      write_address_data_log_force[2793] <= 6'h00;
      write_address_data_log_force[2794] <= 6'h00;
      write_address_data_log_force[2795] <= 6'h00;
      write_address_data_log_force[2796] <= 6'h00;
      write_address_data_log_force[2797] <= 6'h00;
      write_address_data_log_force[2798] <= 6'h00;
      write_address_data_log_force[2799] <= 6'h00;
      write_address_data_log_force[2800] <= 6'h00;
      write_address_data_log_force[2801] <= 6'h00;
      write_address_data_log_force[2802] <= 6'h00;
      write_address_data_log_force[2803] <= 6'h00;
      write_address_data_log_force[2804] <= 6'h00;
      write_address_data_log_force[2805] <= 6'h00;
      write_address_data_log_force[2806] <= 6'h00;
      write_address_data_log_force[2807] <= 6'h00;
      write_address_data_log_force[2808] <= 6'h00;
      write_address_data_log_force[2809] <= 6'h00;
      write_address_data_log_force[2810] <= 6'h00;
      write_address_data_log_force[2811] <= 6'h00;
      write_address_data_log_force[2812] <= 6'h00;
      write_address_data_log_force[2813] <= 6'h00;
      write_address_data_log_force[2814] <= 6'h00;
      write_address_data_log_force[2815] <= 6'h00;
      write_address_data_log_force[2816] <= 6'h00;
      write_address_data_log_force[2817] <= 6'h00;
      write_address_data_log_force[2818] <= 6'h00;
      write_address_data_log_force[2819] <= 6'h00;
      write_address_data_log_force[2820] <= 6'h00;
      write_address_data_log_force[2821] <= 6'h00;
      write_address_data_log_force[2822] <= 6'h00;
      write_address_data_log_force[2823] <= 6'h00;
      write_address_data_log_force[2824] <= 6'h00;
      write_address_data_log_force[2825] <= 6'h00;
      write_address_data_log_force[2826] <= 6'h00;
      write_address_data_log_force[2827] <= 6'h00;
      write_address_data_log_force[2828] <= 6'h00;
      write_address_data_log_force[2829] <= 6'h00;
      write_address_data_log_force[2830] <= 6'h00;
      write_address_data_log_force[2831] <= 6'h00;
      write_address_data_log_force[2832] <= 6'h00;
      write_address_data_log_force[2833] <= 6'h00;
      write_address_data_log_force[2834] <= 6'h00;
      write_address_data_log_force[2835] <= 6'h00;
      write_address_data_log_force[2836] <= 6'h00;
      write_address_data_log_force[2837] <= 6'h00;
      write_address_data_log_force[2838] <= 6'h00;
      write_address_data_log_force[2839] <= 6'h00;
      write_address_data_log_force[2840] <= 6'h00;
      write_address_data_log_force[2841] <= 6'h00;
      write_address_data_log_force[2842] <= 6'h00;
      write_address_data_log_force[2843] <= 6'h00;
      write_address_data_log_force[2844] <= 6'h00;
      write_address_data_log_force[2845] <= 6'h00;
      write_address_data_log_force[2846] <= 6'h00;
      write_address_data_log_force[2847] <= 6'h00;
      write_address_data_log_force[2848] <= 6'h00;
      write_address_data_log_force[2849] <= 6'h00;
      write_address_data_log_force[2850] <= 6'h00;
      write_address_data_log_force[2851] <= 6'h00;
      write_address_data_log_force[2852] <= 6'h00;
      write_address_data_log_force[2853] <= 6'h00;
      write_address_data_log_force[2854] <= 6'h00;
      write_address_data_log_force[2855] <= 6'h00;
      write_address_data_log_force[2856] <= 6'h00;
      write_address_data_log_force[2857] <= 6'h00;
      write_address_data_log_force[2858] <= 6'h00;
      write_address_data_log_force[2859] <= 6'h00;
      write_address_data_log_force[2860] <= 6'h00;
      write_address_data_log_force[2861] <= 6'h00;
      write_address_data_log_force[2862] <= 6'h00;
      write_address_data_log_force[2863] <= 6'h00;
      write_address_data_log_force[2864] <= 6'h00;
      write_address_data_log_force[2865] <= 6'h00;
      write_address_data_log_force[2866] <= 6'h00;
      write_address_data_log_force[2867] <= 6'h00;
      write_address_data_log_force[2868] <= 6'h00;
      write_address_data_log_force[2869] <= 6'h00;
      write_address_data_log_force[2870] <= 6'h00;
      write_address_data_log_force[2871] <= 6'h00;
      write_address_data_log_force[2872] <= 6'h00;
      write_address_data_log_force[2873] <= 6'h00;
      write_address_data_log_force[2874] <= 6'h00;
      write_address_data_log_force[2875] <= 6'h00;
      write_address_data_log_force[2876] <= 6'h00;
      write_address_data_log_force[2877] <= 6'h00;
      write_address_data_log_force[2878] <= 6'h00;
      write_address_data_log_force[2879] <= 6'h00;
      write_address_data_log_force[2880] <= 6'h00;
      write_address_data_log_force[2881] <= 6'h00;
      write_address_data_log_force[2882] <= 6'h00;
      write_address_data_log_force[2883] <= 6'h00;
      write_address_data_log_force[2884] <= 6'h00;
      write_address_data_log_force[2885] <= 6'h00;
      write_address_data_log_force[2886] <= 6'h00;
      write_address_data_log_force[2887] <= 6'h00;
      write_address_data_log_force[2888] <= 6'h00;
      write_address_data_log_force[2889] <= 6'h00;
      write_address_data_log_force[2890] <= 6'h00;
      write_address_data_log_force[2891] <= 6'h00;
      write_address_data_log_force[2892] <= 6'h00;
      write_address_data_log_force[2893] <= 6'h00;
      write_address_data_log_force[2894] <= 6'h00;
      write_address_data_log_force[2895] <= 6'h00;
      write_address_data_log_force[2896] <= 6'h00;
      write_address_data_log_force[2897] <= 6'h00;
      write_address_data_log_force[2898] <= 6'h00;
      write_address_data_log_force[2899] <= 6'h00;
      write_address_data_log_force[2900] <= 6'h00;
      write_address_data_log_force[2901] <= 6'h00;
      write_address_data_log_force[2902] <= 6'h00;
      write_address_data_log_force[2903] <= 6'h00;
      write_address_data_log_force[2904] <= 6'h00;
      write_address_data_log_force[2905] <= 6'h00;
      write_address_data_log_force[2906] <= 6'h00;
      write_address_data_log_force[2907] <= 6'h00;
      write_address_data_log_force[2908] <= 6'h00;
      write_address_data_log_force[2909] <= 6'h00;
      write_address_data_log_force[2910] <= 6'h00;
      write_address_data_log_force[2911] <= 6'h00;
      write_address_data_log_force[2912] <= 6'h00;
      write_address_data_log_force[2913] <= 6'h00;
      write_address_data_log_force[2914] <= 6'h00;
      write_address_data_log_force[2915] <= 6'h00;
      write_address_data_log_force[2916] <= 6'h00;
      write_address_data_log_force[2917] <= 6'h00;
      write_address_data_log_force[2918] <= 6'h00;
      write_address_data_log_force[2919] <= 6'h00;
      write_address_data_log_force[2920] <= 6'h00;
      write_address_data_log_force[2921] <= 6'h00;
      write_address_data_log_force[2922] <= 6'h00;
      write_address_data_log_force[2923] <= 6'h00;
      write_address_data_log_force[2924] <= 6'h00;
      write_address_data_log_force[2925] <= 6'h00;
      write_address_data_log_force[2926] <= 6'h00;
      write_address_data_log_force[2927] <= 6'h00;
      write_address_data_log_force[2928] <= 6'h00;
      write_address_data_log_force[2929] <= 6'h00;
      write_address_data_log_force[2930] <= 6'h00;
      write_address_data_log_force[2931] <= 6'h00;
      write_address_data_log_force[2932] <= 6'h00;
      write_address_data_log_force[2933] <= 6'h00;
      write_address_data_log_force[2934] <= 6'h00;
      write_address_data_log_force[2935] <= 6'h00;
      write_address_data_log_force[2936] <= 6'h00;
      write_address_data_log_force[2937] <= 6'h00;
      write_address_data_log_force[2938] <= 6'h00;
      write_address_data_log_force[2939] <= 6'h00;
      write_address_data_log_force[2940] <= 6'h00;
      write_address_data_log_force[2941] <= 6'h00;
      write_address_data_log_force[2942] <= 6'h00;
      write_address_data_log_force[2943] <= 6'h00;
      write_address_data_log_force[2944] <= 6'h00;
      write_address_data_log_force[2945] <= 6'h00;
      write_address_data_log_force[2946] <= 6'h00;
      write_address_data_log_force[2947] <= 6'h00;
      write_address_data_log_force[2948] <= 6'h00;
      write_address_data_log_force[2949] <= 6'h00;
      write_address_data_log_force[2950] <= 6'h00;
      write_address_data_log_force[2951] <= 6'h00;
      write_address_data_log_force[2952] <= 6'h00;
      write_address_data_log_force[2953] <= 6'h00;
      write_address_data_log_force[2954] <= 6'h00;
      write_address_data_log_force[2955] <= 6'h00;
      write_address_data_log_force[2956] <= 6'h00;
      write_address_data_log_force[2957] <= 6'h00;
      write_address_data_log_force[2958] <= 6'h00;
      write_address_data_log_force[2959] <= 6'h00;
      write_address_data_log_force[2960] <= 6'h00;
      write_address_data_log_force[2961] <= 6'h00;
      write_address_data_log_force[2962] <= 6'h00;
      write_address_data_log_force[2963] <= 6'h00;
      write_address_data_log_force[2964] <= 6'h00;
      write_address_data_log_force[2965] <= 6'h00;
      write_address_data_log_force[2966] <= 6'h00;
      write_address_data_log_force[2967] <= 6'h00;
      write_address_data_log_force[2968] <= 6'h00;
      write_address_data_log_force[2969] <= 6'h00;
      write_address_data_log_force[2970] <= 6'h00;
      write_address_data_log_force[2971] <= 6'h00;
      write_address_data_log_force[2972] <= 6'h00;
      write_address_data_log_force[2973] <= 6'h00;
      write_address_data_log_force[2974] <= 6'h00;
      write_address_data_log_force[2975] <= 6'h00;
      write_address_data_log_force[2976] <= 6'h00;
      write_address_data_log_force[2977] <= 6'h00;
      write_address_data_log_force[2978] <= 6'h00;
      write_address_data_log_force[2979] <= 6'h00;
      write_address_data_log_force[2980] <= 6'h00;
      write_address_data_log_force[2981] <= 6'h00;
      write_address_data_log_force[2982] <= 6'h00;
      write_address_data_log_force[2983] <= 6'h00;
      write_address_data_log_force[2984] <= 6'h00;
      write_address_data_log_force[2985] <= 6'h00;
      write_address_data_log_force[2986] <= 6'h00;
      write_address_data_log_force[2987] <= 6'h00;
      write_address_data_log_force[2988] <= 6'h00;
      write_address_data_log_force[2989] <= 6'h00;
      write_address_data_log_force[2990] <= 6'h00;
      write_address_data_log_force[2991] <= 6'h00;
      write_address_data_log_force[2992] <= 6'h00;
      write_address_data_log_force[2993] <= 6'h00;
      write_address_data_log_force[2994] <= 6'h00;
      write_address_data_log_force[2995] <= 6'h00;
      write_address_data_log_force[2996] <= 6'h00;
      write_address_data_log_force[2997] <= 6'h00;
      write_address_data_log_force[2998] <= 6'h00;
      write_address_data_log_force[2999] <= 6'h00;
      write_address_data_log_force[3000] <= 6'h00;
      write_address_data_log_force[3001] <= 6'h00;
      write_address_data_log_force[3002] <= 6'h00;
      write_address_data_log_force[3003] <= 6'h00;
      write_address_data_log_force[3004] <= 6'h00;
      write_address_data_log_force[3005] <= 6'h00;
      write_address_data_log_force[3006] <= 6'h00;
      write_address_data_log_force[3007] <= 6'h00;
      write_address_data_log_force[3008] <= 6'h00;
      write_address_data_log_force[3009] <= 6'h00;
      write_address_data_log_force[3010] <= 6'h00;
      write_address_data_log_force[3011] <= 6'h00;
      write_address_data_log_force[3012] <= 6'h00;
      write_address_data_log_force[3013] <= 6'h00;
      write_address_data_log_force[3014] <= 6'h00;
      write_address_data_log_force[3015] <= 6'h00;
      write_address_data_log_force[3016] <= 6'h00;
      write_address_data_log_force[3017] <= 6'h00;
      write_address_data_log_force[3018] <= 6'h00;
      write_address_data_log_force[3019] <= 6'h00;
      write_address_data_log_force[3020] <= 6'h00;
      write_address_data_log_force[3021] <= 6'h00;
      write_address_data_log_force[3022] <= 6'h00;
      write_address_data_log_force[3023] <= 6'h00;
      write_address_data_log_force[3024] <= 6'h00;
      write_address_data_log_force[3025] <= 6'h00;
      write_address_data_log_force[3026] <= 6'h00;
      write_address_data_log_force[3027] <= 6'h00;
      write_address_data_log_force[3028] <= 6'h00;
      write_address_data_log_force[3029] <= 6'h00;
      write_address_data_log_force[3030] <= 6'h00;
      write_address_data_log_force[3031] <= 6'h00;
      write_address_data_log_force[3032] <= 6'h00;
      write_address_data_log_force[3033] <= 6'h00;
      write_address_data_log_force[3034] <= 6'h00;
      write_address_data_log_force[3035] <= 6'h00;
      write_address_data_log_force[3036] <= 6'h00;
      write_address_data_log_force[3037] <= 6'h00;
      write_address_data_log_force[3038] <= 6'h00;
      write_address_data_log_force[3039] <= 6'h00;
      write_address_data_log_force[3040] <= 6'h00;
      write_address_data_log_force[3041] <= 6'h00;
      write_address_data_log_force[3042] <= 6'h00;
      write_address_data_log_force[3043] <= 6'h00;
      write_address_data_log_force[3044] <= 6'h00;
      write_address_data_log_force[3045] <= 6'h00;
      write_address_data_log_force[3046] <= 6'h00;
      write_address_data_log_force[3047] <= 6'h00;
      write_address_data_log_force[3048] <= 6'h00;
      write_address_data_log_force[3049] <= 6'h00;
      write_address_data_log_force[3050] <= 6'h00;
      write_address_data_log_force[3051] <= 6'h00;
      write_address_data_log_force[3052] <= 6'h00;
      write_address_data_log_force[3053] <= 6'h00;
      write_address_data_log_force[3054] <= 6'h00;
      write_address_data_log_force[3055] <= 6'h00;
      write_address_data_log_force[3056] <= 6'h00;
      write_address_data_log_force[3057] <= 6'h00;
      write_address_data_log_force[3058] <= 6'h00;
      write_address_data_log_force[3059] <= 6'h00;
      write_address_data_log_force[3060] <= 6'h00;
      write_address_data_log_force[3061] <= 6'h00;
      write_address_data_log_force[3062] <= 6'h00;
      write_address_data_log_force[3063] <= 6'h00;
      write_address_data_log_force[3064] <= 6'h00;
      write_address_data_log_force[3065] <= 6'h00;
      write_address_data_log_force[3066] <= 6'h00;
      write_address_data_log_force[3067] <= 6'h00;
      write_address_data_log_force[3068] <= 6'h00;
      write_address_data_log_force[3069] <= 6'h00;
      write_address_data_log_force[3070] <= 6'h00;
      write_address_data_log_force[3071] <= 6'h00;
      write_address_data_log_force[3072] <= 6'h00;
      write_address_data_log_force[3073] <= 6'h00;
      write_address_data_log_force[3074] <= 6'h00;
      write_address_data_log_force[3075] <= 6'h00;
      write_address_data_log_force[3076] <= 6'h00;
      write_address_data_log_force[3077] <= 6'h00;
      write_address_data_log_force[3078] <= 6'h00;
      write_address_data_log_force[3079] <= 6'h00;
      write_address_data_log_force[3080] <= 6'h00;
      write_address_data_log_force[3081] <= 6'h00;
      write_address_data_log_force[3082] <= 6'h00;
      write_address_data_log_force[3083] <= 6'h00;
      write_address_data_log_force[3084] <= 6'h00;
      write_address_data_log_force[3085] <= 6'h00;
      write_address_data_log_force[3086] <= 6'h00;
      write_address_data_log_force[3087] <= 6'h00;
      write_address_data_log_force[3088] <= 6'h00;
      write_address_data_log_force[3089] <= 6'h00;
      write_address_data_log_force[3090] <= 6'h00;
      write_address_data_log_force[3091] <= 6'h00;
      write_address_data_log_force[3092] <= 6'h00;
      write_address_data_log_force[3093] <= 6'h00;
      write_address_data_log_force[3094] <= 6'h00;
      write_address_data_log_force[3095] <= 6'h00;
      write_address_data_log_force[3096] <= 6'h00;
      write_address_data_log_force[3097] <= 6'h00;
      write_address_data_log_force[3098] <= 6'h00;
      write_address_data_log_force[3099] <= 6'h00;
      write_address_data_log_force[3100] <= 6'h00;
      write_address_data_log_force[3101] <= 6'h00;
      write_address_data_log_force[3102] <= 6'h00;
      write_address_data_log_force[3103] <= 6'h00;
      write_address_data_log_force[3104] <= 6'h00;
      write_address_data_log_force[3105] <= 6'h00;
      write_address_data_log_force[3106] <= 6'h00;
      write_address_data_log_force[3107] <= 6'h00;
      write_address_data_log_force[3108] <= 6'h00;
      write_address_data_log_force[3109] <= 6'h00;
      write_address_data_log_force[3110] <= 6'h00;
      write_address_data_log_force[3111] <= 6'h00;
      write_address_data_log_force[3112] <= 6'h00;
      write_address_data_log_force[3113] <= 6'h00;
      write_address_data_log_force[3114] <= 6'h00;
      write_address_data_log_force[3115] <= 6'h00;
      write_address_data_log_force[3116] <= 6'h00;
      write_address_data_log_force[3117] <= 6'h00;
      write_address_data_log_force[3118] <= 6'h00;
      write_address_data_log_force[3119] <= 6'h00;
      write_address_data_log_force[3120] <= 6'h00;
      write_address_data_log_force[3121] <= 6'h00;
      write_address_data_log_force[3122] <= 6'h00;
      write_address_data_log_force[3123] <= 6'h00;
      write_address_data_log_force[3124] <= 6'h00;
      write_address_data_log_force[3125] <= 6'h00;
      write_address_data_log_force[3126] <= 6'h00;
      write_address_data_log_force[3127] <= 6'h00;
      write_address_data_log_force[3128] <= 6'h00;
      write_address_data_log_force[3129] <= 6'h00;
      write_address_data_log_force[3130] <= 6'h00;
      write_address_data_log_force[3131] <= 6'h00;
      write_address_data_log_force[3132] <= 6'h00;
      write_address_data_log_force[3133] <= 6'h00;
      write_address_data_log_force[3134] <= 6'h00;
      write_address_data_log_force[3135] <= 6'h00;
      write_address_data_log_force[3136] <= 6'h00;
      write_address_data_log_force[3137] <= 6'h00;
      write_address_data_log_force[3138] <= 6'h00;
      write_address_data_log_force[3139] <= 6'h00;
      write_address_data_log_force[3140] <= 6'h00;
      write_address_data_log_force[3141] <= 6'h00;
      write_address_data_log_force[3142] <= 6'h00;
      write_address_data_log_force[3143] <= 6'h00;
      write_address_data_log_force[3144] <= 6'h00;
      write_address_data_log_force[3145] <= 6'h00;
      write_address_data_log_force[3146] <= 6'h00;
      write_address_data_log_force[3147] <= 6'h00;
      write_address_data_log_force[3148] <= 6'h00;
      write_address_data_log_force[3149] <= 6'h00;
      write_address_data_log_force[3150] <= 6'h00;
      write_address_data_log_force[3151] <= 6'h00;
      write_address_data_log_force[3152] <= 6'h00;
      write_address_data_log_force[3153] <= 6'h00;
      write_address_data_log_force[3154] <= 6'h00;
      write_address_data_log_force[3155] <= 6'h00;
      write_address_data_log_force[3156] <= 6'h00;
      write_address_data_log_force[3157] <= 6'h00;
      write_address_data_log_force[3158] <= 6'h00;
      write_address_data_log_force[3159] <= 6'h00;
      write_address_data_log_force[3160] <= 6'h00;
      write_address_data_log_force[3161] <= 6'h00;
      write_address_data_log_force[3162] <= 6'h00;
      write_address_data_log_force[3163] <= 6'h00;
      write_address_data_log_force[3164] <= 6'h00;
      write_address_data_log_force[3165] <= 6'h00;
      write_address_data_log_force[3166] <= 6'h00;
      write_address_data_log_force[3167] <= 6'h00;
      write_address_data_log_force[3168] <= 6'h00;
      write_address_data_log_force[3169] <= 6'h00;
      write_address_data_log_force[3170] <= 6'h00;
      write_address_data_log_force[3171] <= 6'h00;
      write_address_data_log_force[3172] <= 6'h00;
      write_address_data_log_force[3173] <= 6'h00;
      write_address_data_log_force[3174] <= 6'h00;
      write_address_data_log_force[3175] <= 6'h00;
      write_address_data_log_force[3176] <= 6'h00;
      write_address_data_log_force[3177] <= 6'h00;
      write_address_data_log_force[3178] <= 6'h00;
      write_address_data_log_force[3179] <= 6'h00;
      write_address_data_log_force[3180] <= 6'h00;
      write_address_data_log_force[3181] <= 6'h00;
      write_address_data_log_force[3182] <= 6'h00;
      write_address_data_log_force[3183] <= 6'h00;
      write_address_data_log_force[3184] <= 6'h00;
      write_address_data_log_force[3185] <= 6'h00;
      write_address_data_log_force[3186] <= 6'h00;
      write_address_data_log_force[3187] <= 6'h00;
      write_address_data_log_force[3188] <= 6'h00;
      write_address_data_log_force[3189] <= 6'h00;
      write_address_data_log_force[3190] <= 6'h00;
      write_address_data_log_force[3191] <= 6'h00;
      write_address_data_log_force[3192] <= 6'h00;
      write_address_data_log_force[3193] <= 6'h00;
      write_address_data_log_force[3194] <= 6'h00;
      write_address_data_log_force[3195] <= 6'h00;
      write_address_data_log_force[3196] <= 6'h00;
      write_address_data_log_force[3197] <= 6'h00;
      write_address_data_log_force[3198] <= 6'h00;
      write_address_data_log_force[3199] <= 6'h00;
      write_address_data_log_force[3200] <= 6'h00;
      write_address_data_log_force[3201] <= 6'h00;
      write_address_data_log_force[3202] <= 6'h00;
      write_address_data_log_force[3203] <= 6'h00;
      write_address_data_log_force[3204] <= 6'h00;
      write_address_data_log_force[3205] <= 6'h00;
      write_address_data_log_force[3206] <= 6'h00;
      write_address_data_log_force[3207] <= 6'h00;
      write_address_data_log_force[3208] <= 6'h00;
      write_address_data_log_force[3209] <= 6'h00;
      write_address_data_log_force[3210] <= 6'h00;
      write_address_data_log_force[3211] <= 6'h00;
      write_address_data_log_force[3212] <= 6'h00;
      write_address_data_log_force[3213] <= 6'h00;
      write_address_data_log_force[3214] <= 6'h00;
      write_address_data_log_force[3215] <= 6'h00;
      write_address_data_log_force[3216] <= 6'h00;
      write_address_data_log_force[3217] <= 6'h00;
      write_address_data_log_force[3218] <= 6'h00;
      write_address_data_log_force[3219] <= 6'h00;
      write_address_data_log_force[3220] <= 6'h00;
      write_address_data_log_force[3221] <= 6'h00;
      write_address_data_log_force[3222] <= 6'h00;
      write_address_data_log_force[3223] <= 6'h00;
      write_address_data_log_force[3224] <= 6'h00;
      write_address_data_log_force[3225] <= 6'h00;
      write_address_data_log_force[3226] <= 6'h00;
      write_address_data_log_force[3227] <= 6'h00;
      write_address_data_log_force[3228] <= 6'h00;
      write_address_data_log_force[3229] <= 6'h00;
      write_address_data_log_force[3230] <= 6'h00;
      write_address_data_log_force[3231] <= 6'h00;
      write_address_data_log_force[3232] <= 6'h00;
      write_address_data_log_force[3233] <= 6'h00;
      write_address_data_log_force[3234] <= 6'h00;
      write_address_data_log_force[3235] <= 6'h00;
      write_address_data_log_force[3236] <= 6'h00;
      write_address_data_log_force[3237] <= 6'h00;
      write_address_data_log_force[3238] <= 6'h00;
      write_address_data_log_force[3239] <= 6'h00;
      write_address_data_log_force[3240] <= 6'h00;
      write_address_data_log_force[3241] <= 6'h00;
      write_address_data_log_force[3242] <= 6'h00;
      write_address_data_log_force[3243] <= 6'h00;
      write_address_data_log_force[3244] <= 6'h00;
      write_address_data_log_force[3245] <= 6'h00;
      write_address_data_log_force[3246] <= 6'h00;
      write_address_data_log_force[3247] <= 6'h00;
      write_address_data_log_force[3248] <= 6'h00;
      write_address_data_log_force[3249] <= 6'h00;
      write_address_data_log_force[3250] <= 6'h00;
      write_address_data_log_force[3251] <= 6'h00;
      write_address_data_log_force[3252] <= 6'h00;
      write_address_data_log_force[3253] <= 6'h00;
      write_address_data_log_force[3254] <= 6'h00;
      write_address_data_log_force[3255] <= 6'h00;
      write_address_data_log_force[3256] <= 6'h00;
      write_address_data_log_force[3257] <= 6'h00;
      write_address_data_log_force[3258] <= 6'h00;
      write_address_data_log_force[3259] <= 6'h00;
      write_address_data_log_force[3260] <= 6'h00;
      write_address_data_log_force[3261] <= 6'h00;
      write_address_data_log_force[3262] <= 6'h00;
      write_address_data_log_force[3263] <= 6'h00;
      write_address_data_log_force[3264] <= 6'h00;
      write_address_data_log_force[3265] <= 6'h00;
      write_address_data_log_force[3266] <= 6'h00;
      write_address_data_log_force[3267] <= 6'h00;
      write_address_data_log_force[3268] <= 6'h00;
      write_address_data_log_force[3269] <= 6'h00;
      write_address_data_log_force[3270] <= 6'h00;
      write_address_data_log_force[3271] <= 6'h00;
      write_address_data_log_force[3272] <= 6'h00;
      write_address_data_log_force[3273] <= 6'h00;
      write_address_data_log_force[3274] <= 6'h00;
      write_address_data_log_force[3275] <= 6'h00;
      write_address_data_log_force[3276] <= 6'h00;
      write_address_data_log_force[3277] <= 6'h00;
      write_address_data_log_force[3278] <= 6'h00;
      write_address_data_log_force[3279] <= 6'h00;
      write_address_data_log_force[3280] <= 6'h00;
      write_address_data_log_force[3281] <= 6'h00;
      write_address_data_log_force[3282] <= 6'h00;
      write_address_data_log_force[3283] <= 6'h00;
      write_address_data_log_force[3284] <= 6'h00;
      write_address_data_log_force[3285] <= 6'h00;
      write_address_data_log_force[3286] <= 6'h00;
      write_address_data_log_force[3287] <= 6'h00;
      write_address_data_log_force[3288] <= 6'h00;
      write_address_data_log_force[3289] <= 6'h00;
      write_address_data_log_force[3290] <= 6'h00;
      write_address_data_log_force[3291] <= 6'h00;
      write_address_data_log_force[3292] <= 6'h00;
      write_address_data_log_force[3293] <= 6'h00;
      write_address_data_log_force[3294] <= 6'h00;
      write_address_data_log_force[3295] <= 6'h00;
      write_address_data_log_force[3296] <= 6'h00;
      write_address_data_log_force[3297] <= 6'h00;
      write_address_data_log_force[3298] <= 6'h00;
      write_address_data_log_force[3299] <= 6'h00;
      write_address_data_log_force[3300] <= 6'h00;
      write_address_data_log_force[3301] <= 6'h00;
      write_address_data_log_force[3302] <= 6'h00;
      write_address_data_log_force[3303] <= 6'h00;
      write_address_data_log_force[3304] <= 6'h00;
      write_address_data_log_force[3305] <= 6'h00;
      write_address_data_log_force[3306] <= 6'h00;
      write_address_data_log_force[3307] <= 6'h00;
      write_address_data_log_force[3308] <= 6'h00;
      write_address_data_log_force[3309] <= 6'h00;
      write_address_data_log_force[3310] <= 6'h00;
      write_address_data_log_force[3311] <= 6'h00;
      write_address_data_log_force[3312] <= 6'h00;
      write_address_data_log_force[3313] <= 6'h00;
      write_address_data_log_force[3314] <= 6'h00;
      write_address_data_log_force[3315] <= 6'h00;
      write_address_data_log_force[3316] <= 6'h00;
      write_address_data_log_force[3317] <= 6'h00;
      write_address_data_log_force[3318] <= 6'h00;
      write_address_data_log_force[3319] <= 6'h00;
      write_address_data_log_force[3320] <= 6'h00;
      write_address_data_log_force[3321] <= 6'h00;
      write_address_data_log_force[3322] <= 6'h00;
      write_address_data_log_force[3323] <= 6'h00;
      write_address_data_log_force[3324] <= 6'h00;
      write_address_data_log_force[3325] <= 6'h00;
      write_address_data_log_force[3326] <= 6'h00;
      write_address_data_log_force[3327] <= 6'h00;
      write_address_data_log_force[3328] <= 6'h00;
      write_address_data_log_force[3329] <= 6'h00;
      write_address_data_log_force[3330] <= 6'h00;
      write_address_data_log_force[3331] <= 6'h00;
      write_address_data_log_force[3332] <= 6'h00;
      write_address_data_log_force[3333] <= 6'h00;
      write_address_data_log_force[3334] <= 6'h00;
      write_address_data_log_force[3335] <= 6'h00;
      write_address_data_log_force[3336] <= 6'h00;
      write_address_data_log_force[3337] <= 6'h00;
      write_address_data_log_force[3338] <= 6'h00;
      write_address_data_log_force[3339] <= 6'h00;
      write_address_data_log_force[3340] <= 6'h00;
      write_address_data_log_force[3341] <= 6'h00;
      write_address_data_log_force[3342] <= 6'h00;
      write_address_data_log_force[3343] <= 6'h00;
      write_address_data_log_force[3344] <= 6'h00;
      write_address_data_log_force[3345] <= 6'h00;
      write_address_data_log_force[3346] <= 6'h00;
      write_address_data_log_force[3347] <= 6'h00;
      write_address_data_log_force[3348] <= 6'h00;
      write_address_data_log_force[3349] <= 6'h00;
      write_address_data_log_force[3350] <= 6'h00;
      write_address_data_log_force[3351] <= 6'h00;
      write_address_data_log_force[3352] <= 6'h00;
      write_address_data_log_force[3353] <= 6'h00;
      write_address_data_log_force[3354] <= 6'h00;
      write_address_data_log_force[3355] <= 6'h00;
      write_address_data_log_force[3356] <= 6'h00;
      write_address_data_log_force[3357] <= 6'h00;
      write_address_data_log_force[3358] <= 6'h00;
      write_address_data_log_force[3359] <= 6'h00;
      write_address_data_log_force[3360] <= 6'h00;
      write_address_data_log_force[3361] <= 6'h00;
      write_address_data_log_force[3362] <= 6'h00;
      write_address_data_log_force[3363] <= 6'h00;
      write_address_data_log_force[3364] <= 6'h00;
      write_address_data_log_force[3365] <= 6'h00;
      write_address_data_log_force[3366] <= 6'h00;
      write_address_data_log_force[3367] <= 6'h00;
      write_address_data_log_force[3368] <= 6'h00;
      write_address_data_log_force[3369] <= 6'h00;
      write_address_data_log_force[3370] <= 6'h00;
      write_address_data_log_force[3371] <= 6'h00;
      write_address_data_log_force[3372] <= 6'h00;
      write_address_data_log_force[3373] <= 6'h00;
      write_address_data_log_force[3374] <= 6'h00;
      write_address_data_log_force[3375] <= 6'h00;
      write_address_data_log_force[3376] <= 6'h00;
      write_address_data_log_force[3377] <= 6'h00;
      write_address_data_log_force[3378] <= 6'h00;
      write_address_data_log_force[3379] <= 6'h00;
      write_address_data_log_force[3380] <= 6'h00;
      write_address_data_log_force[3381] <= 6'h00;
      write_address_data_log_force[3382] <= 6'h00;
      write_address_data_log_force[3383] <= 6'h00;
      write_address_data_log_force[3384] <= 6'h00;
      write_address_data_log_force[3385] <= 6'h00;
      write_address_data_log_force[3386] <= 6'h00;
      write_address_data_log_force[3387] <= 6'h00;
      write_address_data_log_force[3388] <= 6'h00;
      write_address_data_log_force[3389] <= 6'h00;
      write_address_data_log_force[3390] <= 6'h00;
      write_address_data_log_force[3391] <= 6'h00;
      write_address_data_log_force[3392] <= 6'h00;
      write_address_data_log_force[3393] <= 6'h00;
      write_address_data_log_force[3394] <= 6'h00;
      write_address_data_log_force[3395] <= 6'h00;
      write_address_data_log_force[3396] <= 6'h00;
      write_address_data_log_force[3397] <= 6'h00;
      write_address_data_log_force[3398] <= 6'h00;
      write_address_data_log_force[3399] <= 6'h00;
      write_address_data_log_force[3400] <= 6'h00;
      write_address_data_log_force[3401] <= 6'h00;
      write_address_data_log_force[3402] <= 6'h00;
      write_address_data_log_force[3403] <= 6'h00;
      write_address_data_log_force[3404] <= 6'h00;
      write_address_data_log_force[3405] <= 6'h00;
      write_address_data_log_force[3406] <= 6'h00;
      write_address_data_log_force[3407] <= 6'h00;
      write_address_data_log_force[3408] <= 6'h00;
      write_address_data_log_force[3409] <= 6'h00;
      write_address_data_log_force[3410] <= 6'h00;
      write_address_data_log_force[3411] <= 6'h00;
      write_address_data_log_force[3412] <= 6'h00;
      write_address_data_log_force[3413] <= 6'h00;
      write_address_data_log_force[3414] <= 6'h00;
      write_address_data_log_force[3415] <= 6'h00;
      write_address_data_log_force[3416] <= 6'h00;
      write_address_data_log_force[3417] <= 6'h00;
      write_address_data_log_force[3418] <= 6'h00;
      write_address_data_log_force[3419] <= 6'h00;
      write_address_data_log_force[3420] <= 6'h00;
      write_address_data_log_force[3421] <= 6'h00;
      write_address_data_log_force[3422] <= 6'h00;
      write_address_data_log_force[3423] <= 6'h00;
      write_address_data_log_force[3424] <= 6'h00;
      write_address_data_log_force[3425] <= 6'h00;
      write_address_data_log_force[3426] <= 6'h00;
      write_address_data_log_force[3427] <= 6'h00;
      write_address_data_log_force[3428] <= 6'h00;
      write_address_data_log_force[3429] <= 6'h00;
      write_address_data_log_force[3430] <= 6'h00;
      write_address_data_log_force[3431] <= 6'h00;
      write_address_data_log_force[3432] <= 6'h00;
      write_address_data_log_force[3433] <= 6'h00;
      write_address_data_log_force[3434] <= 6'h00;
      write_address_data_log_force[3435] <= 6'h00;
      write_address_data_log_force[3436] <= 6'h00;
      write_address_data_log_force[3437] <= 6'h00;
      write_address_data_log_force[3438] <= 6'h00;
      write_address_data_log_force[3439] <= 6'h00;
      write_address_data_log_force[3440] <= 6'h00;
      write_address_data_log_force[3441] <= 6'h00;
      write_address_data_log_force[3442] <= 6'h00;
      write_address_data_log_force[3443] <= 6'h00;
      write_address_data_log_force[3444] <= 6'h00;
      write_address_data_log_force[3445] <= 6'h00;
      write_address_data_log_force[3446] <= 6'h00;
      write_address_data_log_force[3447] <= 6'h00;
      write_address_data_log_force[3448] <= 6'h00;
      write_address_data_log_force[3449] <= 6'h00;
      write_address_data_log_force[3450] <= 6'h00;
      write_address_data_log_force[3451] <= 6'h00;
      write_address_data_log_force[3452] <= 6'h00;
      write_address_data_log_force[3453] <= 6'h00;
      write_address_data_log_force[3454] <= 6'h00;
      write_address_data_log_force[3455] <= 6'h00;
      write_address_data_log_force[3456] <= 6'h00;
      write_address_data_log_force[3457] <= 6'h00;
      write_address_data_log_force[3458] <= 6'h00;
      write_address_data_log_force[3459] <= 6'h00;
      write_address_data_log_force[3460] <= 6'h00;
      write_address_data_log_force[3461] <= 6'h00;
      write_address_data_log_force[3462] <= 6'h00;
      write_address_data_log_force[3463] <= 6'h00;
      write_address_data_log_force[3464] <= 6'h00;
      write_address_data_log_force[3465] <= 6'h00;
      write_address_data_log_force[3466] <= 6'h00;
      write_address_data_log_force[3467] <= 6'h00;
      write_address_data_log_force[3468] <= 6'h00;
      write_address_data_log_force[3469] <= 6'h00;
      write_address_data_log_force[3470] <= 6'h00;
      write_address_data_log_force[3471] <= 6'h00;
      write_address_data_log_force[3472] <= 6'h00;
      write_address_data_log_force[3473] <= 6'h00;
      write_address_data_log_force[3474] <= 6'h00;
      write_address_data_log_force[3475] <= 6'h00;
      write_address_data_log_force[3476] <= 6'h00;
      write_address_data_log_force[3477] <= 6'h00;
      write_address_data_log_force[3478] <= 6'h00;
      write_address_data_log_force[3479] <= 6'h00;
      write_address_data_log_force[3480] <= 6'h00;
      write_address_data_log_force[3481] <= 6'h00;
      write_address_data_log_force[3482] <= 6'h00;
      write_address_data_log_force[3483] <= 6'h00;
      write_address_data_log_force[3484] <= 6'h00;
      write_address_data_log_force[3485] <= 6'h00;
      write_address_data_log_force[3486] <= 6'h00;
      write_address_data_log_force[3487] <= 6'h00;
      write_address_data_log_force[3488] <= 6'h00;
      write_address_data_log_force[3489] <= 6'h00;
      write_address_data_log_force[3490] <= 6'h00;
      write_address_data_log_force[3491] <= 6'h00;
      write_address_data_log_force[3492] <= 6'h00;
      write_address_data_log_force[3493] <= 6'h00;
      write_address_data_log_force[3494] <= 6'h00;
      write_address_data_log_force[3495] <= 6'h00;
      write_address_data_log_force[3496] <= 6'h00;
      write_address_data_log_force[3497] <= 6'h00;
      write_address_data_log_force[3498] <= 6'h00;
      write_address_data_log_force[3499] <= 6'h00;
      write_address_data_log_force[3500] <= 6'h00;
      write_address_data_log_force[3501] <= 6'h00;
      write_address_data_log_force[3502] <= 6'h00;
      write_address_data_log_force[3503] <= 6'h00;
      write_address_data_log_force[3504] <= 6'h00;
      write_address_data_log_force[3505] <= 6'h00;
      write_address_data_log_force[3506] <= 6'h00;
      write_address_data_log_force[3507] <= 6'h00;
      write_address_data_log_force[3508] <= 6'h00;
      write_address_data_log_force[3509] <= 6'h00;
      write_address_data_log_force[3510] <= 6'h00;
      write_address_data_log_force[3511] <= 6'h00;
      write_address_data_log_force[3512] <= 6'h00;
      write_address_data_log_force[3513] <= 6'h00;
      write_address_data_log_force[3514] <= 6'h00;
      write_address_data_log_force[3515] <= 6'h00;
      write_address_data_log_force[3516] <= 6'h00;
      write_address_data_log_force[3517] <= 6'h00;
      write_address_data_log_force[3518] <= 6'h00;
      write_address_data_log_force[3519] <= 6'h00;
      write_address_data_log_force[3520] <= 6'h00;
      write_address_data_log_force[3521] <= 6'h00;
      write_address_data_log_force[3522] <= 6'h00;
      write_address_data_log_force[3523] <= 6'h00;
      write_address_data_log_force[3524] <= 6'h00;
      write_address_data_log_force[3525] <= 6'h00;
      write_address_data_log_force[3526] <= 6'h00;
      write_address_data_log_force[3527] <= 6'h00;
      write_address_data_log_force[3528] <= 6'h00;
      write_address_data_log_force[3529] <= 6'h00;
      write_address_data_log_force[3530] <= 6'h00;
      write_address_data_log_force[3531] <= 6'h00;
      write_address_data_log_force[3532] <= 6'h00;
      write_address_data_log_force[3533] <= 6'h00;
      write_address_data_log_force[3534] <= 6'h00;
      write_address_data_log_force[3535] <= 6'h00;
      write_address_data_log_force[3536] <= 6'h00;
      write_address_data_log_force[3537] <= 6'h00;
      write_address_data_log_force[3538] <= 6'h00;
      write_address_data_log_force[3539] <= 6'h00;
      write_address_data_log_force[3540] <= 6'h00;
      write_address_data_log_force[3541] <= 6'h00;
      write_address_data_log_force[3542] <= 6'h00;
      write_address_data_log_force[3543] <= 6'h00;
      write_address_data_log_force[3544] <= 6'h00;
      write_address_data_log_force[3545] <= 6'h00;
      write_address_data_log_force[3546] <= 6'h00;
      write_address_data_log_force[3547] <= 6'h00;
      write_address_data_log_force[3548] <= 6'h00;
      write_address_data_log_force[3549] <= 6'h00;
      write_address_data_log_force[3550] <= 6'h00;
      write_address_data_log_force[3551] <= 6'h00;
      write_address_data_log_force[3552] <= 6'h00;
      write_address_data_log_force[3553] <= 6'h00;
      write_address_data_log_force[3554] <= 6'h00;
      write_address_data_log_force[3555] <= 6'h00;
      write_address_data_log_force[3556] <= 6'h00;
      write_address_data_log_force[3557] <= 6'h00;
      write_address_data_log_force[3558] <= 6'h00;
      write_address_data_log_force[3559] <= 6'h00;
      write_address_data_log_force[3560] <= 6'h00;
      write_address_data_log_force[3561] <= 6'h00;
      write_address_data_log_force[3562] <= 6'h00;
      write_address_data_log_force[3563] <= 6'h00;
      write_address_data_log_force[3564] <= 6'h00;
      write_address_data_log_force[3565] <= 6'h00;
      write_address_data_log_force[3566] <= 6'h00;
      write_address_data_log_force[3567] <= 6'h00;
      write_address_data_log_force[3568] <= 6'h00;
      write_address_data_log_force[3569] <= 6'h00;
      write_address_data_log_force[3570] <= 6'h00;
      write_address_data_log_force[3571] <= 6'h00;
      write_address_data_log_force[3572] <= 6'h00;
      write_address_data_log_force[3573] <= 6'h00;
      write_address_data_log_force[3574] <= 6'h00;
      write_address_data_log_force[3575] <= 6'h00;
      write_address_data_log_force[3576] <= 6'h00;
      write_address_data_log_force[3577] <= 6'h00;
      write_address_data_log_force[3578] <= 6'h00;
      write_address_data_log_force[3579] <= 6'h00;
      write_address_data_log_force[3580] <= 6'h00;
      write_address_data_log_force[3581] <= 6'h00;
      write_address_data_log_force[3582] <= 6'h00;
      write_address_data_log_force[3583] <= 6'h00;
      write_address_data_log_force[3584] <= 6'h00;
      write_address_data_log_force[3585] <= 6'h00;
      write_address_data_log_force[3586] <= 6'h00;
      write_address_data_log_force[3587] <= 6'h00;
      write_address_data_log_force[3588] <= 6'h00;
      write_address_data_log_force[3589] <= 6'h00;
      write_address_data_log_force[3590] <= 6'h00;
      write_address_data_log_force[3591] <= 6'h00;
      write_address_data_log_force[3592] <= 6'h00;
      write_address_data_log_force[3593] <= 6'h00;
      write_address_data_log_force[3594] <= 6'h00;
      write_address_data_log_force[3595] <= 6'h00;
      write_address_data_log_force[3596] <= 6'h00;
      write_address_data_log_force[3597] <= 6'h00;
      write_address_data_log_force[3598] <= 6'h00;
      write_address_data_log_force[3599] <= 6'h00;
      write_address_data_log_force[3600] <= 6'h00;
      write_address_data_log_force[3601] <= 6'h00;
      write_address_data_log_force[3602] <= 6'h00;
      write_address_data_log_force[3603] <= 6'h00;
      write_address_data_log_force[3604] <= 6'h00;
      write_address_data_log_force[3605] <= 6'h00;
      write_address_data_log_force[3606] <= 6'h00;
      write_address_data_log_force[3607] <= 6'h00;
      write_address_data_log_force[3608] <= 6'h00;
      write_address_data_log_force[3609] <= 6'h00;
      write_address_data_log_force[3610] <= 6'h00;
      write_address_data_log_force[3611] <= 6'h00;
      write_address_data_log_force[3612] <= 6'h00;
      write_address_data_log_force[3613] <= 6'h00;
      write_address_data_log_force[3614] <= 6'h00;
      write_address_data_log_force[3615] <= 6'h00;
      write_address_data_log_force[3616] <= 6'h00;
      write_address_data_log_force[3617] <= 6'h00;
      write_address_data_log_force[3618] <= 6'h00;
      write_address_data_log_force[3619] <= 6'h00;
      write_address_data_log_force[3620] <= 6'h00;
      write_address_data_log_force[3621] <= 6'h00;
      write_address_data_log_force[3622] <= 6'h00;
      write_address_data_log_force[3623] <= 6'h00;
      write_address_data_log_force[3624] <= 6'h00;
      write_address_data_log_force[3625] <= 6'h00;
      write_address_data_log_force[3626] <= 6'h00;
      write_address_data_log_force[3627] <= 6'h00;
      write_address_data_log_force[3628] <= 6'h00;
      write_address_data_log_force[3629] <= 6'h00;
      write_address_data_log_force[3630] <= 6'h00;
      write_address_data_log_force[3631] <= 6'h00;
      write_address_data_log_force[3632] <= 6'h00;
      write_address_data_log_force[3633] <= 6'h00;
      write_address_data_log_force[3634] <= 6'h00;
      write_address_data_log_force[3635] <= 6'h00;
      write_address_data_log_force[3636] <= 6'h00;
      write_address_data_log_force[3637] <= 6'h00;
      write_address_data_log_force[3638] <= 6'h00;
      write_address_data_log_force[3639] <= 6'h00;
      write_address_data_log_force[3640] <= 6'h00;
      write_address_data_log_force[3641] <= 6'h00;
      write_address_data_log_force[3642] <= 6'h00;
      write_address_data_log_force[3643] <= 6'h00;
      write_address_data_log_force[3644] <= 6'h00;
      write_address_data_log_force[3645] <= 6'h00;
      write_address_data_log_force[3646] <= 6'h00;
      write_address_data_log_force[3647] <= 6'h00;
      write_address_data_log_force[3648] <= 6'h00;
      write_address_data_log_force[3649] <= 6'h00;
      write_address_data_log_force[3650] <= 6'h00;
      write_address_data_log_force[3651] <= 6'h00;
      write_address_data_log_force[3652] <= 6'h00;
      write_address_data_log_force[3653] <= 6'h00;
      write_address_data_log_force[3654] <= 6'h00;
      write_address_data_log_force[3655] <= 6'h00;
      write_address_data_log_force[3656] <= 6'h00;
      write_address_data_log_force[3657] <= 6'h00;
      write_address_data_log_force[3658] <= 6'h00;
      write_address_data_log_force[3659] <= 6'h00;
      write_address_data_log_force[3660] <= 6'h00;
      write_address_data_log_force[3661] <= 6'h00;
      write_address_data_log_force[3662] <= 6'h00;
      write_address_data_log_force[3663] <= 6'h00;
      write_address_data_log_force[3664] <= 6'h00;
      write_address_data_log_force[3665] <= 6'h00;
      write_address_data_log_force[3666] <= 6'h00;
      write_address_data_log_force[3667] <= 6'h00;
      write_address_data_log_force[3668] <= 6'h00;
      write_address_data_log_force[3669] <= 6'h00;
      write_address_data_log_force[3670] <= 6'h00;
      write_address_data_log_force[3671] <= 6'h00;
      write_address_data_log_force[3672] <= 6'h00;
      write_address_data_log_force[3673] <= 6'h00;
      write_address_data_log_force[3674] <= 6'h00;
      write_address_data_log_force[3675] <= 6'h00;
      write_address_data_log_force[3676] <= 6'h00;
      write_address_data_log_force[3677] <= 6'h00;
      write_address_data_log_force[3678] <= 6'h00;
      write_address_data_log_force[3679] <= 6'h00;
      write_address_data_log_force[3680] <= 6'h00;
      write_address_data_log_force[3681] <= 6'h00;
      write_address_data_log_force[3682] <= 6'h00;
      write_address_data_log_force[3683] <= 6'h00;
      write_address_data_log_force[3684] <= 6'h00;
      write_address_data_log_force[3685] <= 6'h00;
      write_address_data_log_force[3686] <= 6'h00;
      write_address_data_log_force[3687] <= 6'h00;
      write_address_data_log_force[3688] <= 6'h00;
      write_address_data_log_force[3689] <= 6'h00;
      write_address_data_log_force[3690] <= 6'h00;
      write_address_data_log_force[3691] <= 6'h00;
      write_address_data_log_force[3692] <= 6'h00;
      write_address_data_log_force[3693] <= 6'h00;
      write_address_data_log_force[3694] <= 6'h00;
      write_address_data_log_force[3695] <= 6'h00;
      write_address_data_log_force[3696] <= 6'h00;
      write_address_data_log_force[3697] <= 6'h00;
      write_address_data_log_force[3698] <= 6'h00;
      write_address_data_log_force[3699] <= 6'h00;
      write_address_data_log_force[3700] <= 6'h00;
      write_address_data_log_force[3701] <= 6'h00;
      write_address_data_log_force[3702] <= 6'h00;
      write_address_data_log_force[3703] <= 6'h00;
      write_address_data_log_force[3704] <= 6'h00;
      write_address_data_log_force[3705] <= 6'h00;
      write_address_data_log_force[3706] <= 6'h00;
      write_address_data_log_force[3707] <= 6'h00;
      write_address_data_log_force[3708] <= 6'h00;
      write_address_data_log_force[3709] <= 6'h00;
      write_address_data_log_force[3710] <= 6'h00;
      write_address_data_log_force[3711] <= 6'h00;
      write_address_data_log_force[3712] <= 6'h00;
      write_address_data_log_force[3713] <= 6'h00;
      write_address_data_log_force[3714] <= 6'h00;
      write_address_data_log_force[3715] <= 6'h00;
      write_address_data_log_force[3716] <= 6'h00;
      write_address_data_log_force[3717] <= 6'h00;
      write_address_data_log_force[3718] <= 6'h00;
      write_address_data_log_force[3719] <= 6'h00;
      write_address_data_log_force[3720] <= 6'h00;
      write_address_data_log_force[3721] <= 6'h00;
      write_address_data_log_force[3722] <= 6'h00;
      write_address_data_log_force[3723] <= 6'h00;
      write_address_data_log_force[3724] <= 6'h00;
      write_address_data_log_force[3725] <= 6'h00;
      write_address_data_log_force[3726] <= 6'h00;
      write_address_data_log_force[3727] <= 6'h00;
      write_address_data_log_force[3728] <= 6'h00;
      write_address_data_log_force[3729] <= 6'h00;
      write_address_data_log_force[3730] <= 6'h00;
      write_address_data_log_force[3731] <= 6'h00;
      write_address_data_log_force[3732] <= 6'h00;
      write_address_data_log_force[3733] <= 6'h00;
      write_address_data_log_force[3734] <= 6'h00;
      write_address_data_log_force[3735] <= 6'h00;
      write_address_data_log_force[3736] <= 6'h00;
      write_address_data_log_force[3737] <= 6'h00;
      write_address_data_log_force[3738] <= 6'h00;
      write_address_data_log_force[3739] <= 6'h00;
      write_address_data_log_force[3740] <= 6'h00;
      write_address_data_log_force[3741] <= 6'h00;
      write_address_data_log_force[3742] <= 6'h00;
      write_address_data_log_force[3743] <= 6'h00;
      write_address_data_log_force[3744] <= 6'h00;
      write_address_data_log_force[3745] <= 6'h00;
      write_address_data_log_force[3746] <= 6'h00;
      write_address_data_log_force[3747] <= 6'h00;
      write_address_data_log_force[3748] <= 6'h00;
      write_address_data_log_force[3749] <= 6'h00;
      write_address_data_log_force[3750] <= 6'h00;
      write_address_data_log_force[3751] <= 6'h00;
      write_address_data_log_force[3752] <= 6'h00;
      write_address_data_log_force[3753] <= 6'h00;
      write_address_data_log_force[3754] <= 6'h00;
      write_address_data_log_force[3755] <= 6'h00;
      write_address_data_log_force[3756] <= 6'h00;
      write_address_data_log_force[3757] <= 6'h00;
      write_address_data_log_force[3758] <= 6'h00;
      write_address_data_log_force[3759] <= 6'h00;
      write_address_data_log_force[3760] <= 6'h00;
      write_address_data_log_force[3761] <= 6'h00;
      write_address_data_log_force[3762] <= 6'h00;
      write_address_data_log_force[3763] <= 6'h00;
      write_address_data_log_force[3764] <= 6'h00;
      write_address_data_log_force[3765] <= 6'h00;
      write_address_data_log_force[3766] <= 6'h00;
      write_address_data_log_force[3767] <= 6'h00;
      write_address_data_log_force[3768] <= 6'h00;
      write_address_data_log_force[3769] <= 6'h00;
      write_address_data_log_force[3770] <= 6'h00;
      write_address_data_log_force[3771] <= 6'h00;
      write_address_data_log_force[3772] <= 6'h00;
      write_address_data_log_force[3773] <= 6'h00;
      write_address_data_log_force[3774] <= 6'h00;
      write_address_data_log_force[3775] <= 6'h00;
      write_address_data_log_force[3776] <= 6'h00;
      write_address_data_log_force[3777] <= 6'h00;
      write_address_data_log_force[3778] <= 6'h00;
      write_address_data_log_force[3779] <= 6'h00;
      write_address_data_log_force[3780] <= 6'h00;
      write_address_data_log_force[3781] <= 6'h00;
      write_address_data_log_force[3782] <= 6'h00;
      write_address_data_log_force[3783] <= 6'h00;
      write_address_data_log_force[3784] <= 6'h00;
      write_address_data_log_force[3785] <= 6'h00;
      write_address_data_log_force[3786] <= 6'h00;
      write_address_data_log_force[3787] <= 6'h00;
      write_address_data_log_force[3788] <= 6'h00;
      write_address_data_log_force[3789] <= 6'h00;
      write_address_data_log_force[3790] <= 6'h00;
      write_address_data_log_force[3791] <= 6'h00;
      write_address_data_log_force[3792] <= 6'h00;
      write_address_data_log_force[3793] <= 6'h00;
      write_address_data_log_force[3794] <= 6'h00;
      write_address_data_log_force[3795] <= 6'h00;
      write_address_data_log_force[3796] <= 6'h00;
      write_address_data_log_force[3797] <= 6'h00;
      write_address_data_log_force[3798] <= 6'h00;
      write_address_data_log_force[3799] <= 6'h00;
      write_address_data_log_force[3800] <= 6'h00;
      write_address_data_log_force[3801] <= 6'h00;
      write_address_data_log_force[3802] <= 6'h00;
      write_address_data_log_force[3803] <= 6'h00;
      write_address_data_log_force[3804] <= 6'h00;
      write_address_data_log_force[3805] <= 6'h00;
      write_address_data_log_force[3806] <= 6'h00;
      write_address_data_log_force[3807] <= 6'h00;
      write_address_data_log_force[3808] <= 6'h00;
      write_address_data_log_force[3809] <= 6'h00;
      write_address_data_log_force[3810] <= 6'h00;
      write_address_data_log_force[3811] <= 6'h00;
      write_address_data_log_force[3812] <= 6'h00;
      write_address_data_log_force[3813] <= 6'h00;
      write_address_data_log_force[3814] <= 6'h00;
      write_address_data_log_force[3815] <= 6'h00;
      write_address_data_log_force[3816] <= 6'h00;
      write_address_data_log_force[3817] <= 6'h00;
      write_address_data_log_force[3818] <= 6'h00;
      write_address_data_log_force[3819] <= 6'h00;
      write_address_data_log_force[3820] <= 6'h00;
      write_address_data_log_force[3821] <= 6'h00;
      write_address_data_log_force[3822] <= 6'h00;
      write_address_data_log_force[3823] <= 6'h00;
      write_address_data_log_force[3824] <= 6'h00;
      write_address_data_log_force[3825] <= 6'h00;
      write_address_data_log_force[3826] <= 6'h00;
      write_address_data_log_force[3827] <= 6'h00;
      write_address_data_log_force[3828] <= 6'h00;
      write_address_data_log_force[3829] <= 6'h00;
      write_address_data_log_force[3830] <= 6'h00;
      write_address_data_log_force[3831] <= 6'h00;
      write_address_data_log_force[3832] <= 6'h00;
      write_address_data_log_force[3833] <= 6'h00;
      write_address_data_log_force[3834] <= 6'h00;
      write_address_data_log_force[3835] <= 6'h00;
      write_address_data_log_force[3836] <= 6'h00;
      write_address_data_log_force[3837] <= 6'h00;
      write_address_data_log_force[3838] <= 6'h00;
      write_address_data_log_force[3839] <= 6'h00;
      write_address_data_log_force[3840] <= 6'h00;
      write_address_data_log_force[3841] <= 6'h00;
      write_address_data_log_force[3842] <= 6'h00;
      write_address_data_log_force[3843] <= 6'h00;
      write_address_data_log_force[3844] <= 6'h00;
      write_address_data_log_force[3845] <= 6'h00;
      write_address_data_log_force[3846] <= 6'h00;
      write_address_data_log_force[3847] <= 6'h00;
      write_address_data_log_force[3848] <= 6'h00;
      write_address_data_log_force[3849] <= 6'h00;
      write_address_data_log_force[3850] <= 6'h00;
      write_address_data_log_force[3851] <= 6'h00;
      write_address_data_log_force[3852] <= 6'h00;
      write_address_data_log_force[3853] <= 6'h00;
      write_address_data_log_force[3854] <= 6'h00;
      write_address_data_log_force[3855] <= 6'h00;
      write_address_data_log_force[3856] <= 6'h00;
      write_address_data_log_force[3857] <= 6'h00;
      write_address_data_log_force[3858] <= 6'h00;
      write_address_data_log_force[3859] <= 6'h00;
      write_address_data_log_force[3860] <= 6'h00;
      write_address_data_log_force[3861] <= 6'h00;
      write_address_data_log_force[3862] <= 6'h00;
      write_address_data_log_force[3863] <= 6'h00;
      write_address_data_log_force[3864] <= 6'h00;
      write_address_data_log_force[3865] <= 6'h00;
      write_address_data_log_force[3866] <= 6'h00;
      write_address_data_log_force[3867] <= 6'h00;
      write_address_data_log_force[3868] <= 6'h00;
      write_address_data_log_force[3869] <= 6'h00;
      write_address_data_log_force[3870] <= 6'h00;
      write_address_data_log_force[3871] <= 6'h00;
      write_address_data_log_force[3872] <= 6'h00;
      write_address_data_log_force[3873] <= 6'h00;
      write_address_data_log_force[3874] <= 6'h00;
      write_address_data_log_force[3875] <= 6'h00;
      write_address_data_log_force[3876] <= 6'h00;
      write_address_data_log_force[3877] <= 6'h00;
      write_address_data_log_force[3878] <= 6'h00;
      write_address_data_log_force[3879] <= 6'h00;
      write_address_data_log_force[3880] <= 6'h00;
      write_address_data_log_force[3881] <= 6'h00;
      write_address_data_log_force[3882] <= 6'h00;
      write_address_data_log_force[3883] <= 6'h00;
      write_address_data_log_force[3884] <= 6'h00;
      write_address_data_log_force[3885] <= 6'h00;
      write_address_data_log_force[3886] <= 6'h00;
      write_address_data_log_force[3887] <= 6'h00;
      write_address_data_log_force[3888] <= 6'h00;
      write_address_data_log_force[3889] <= 6'h00;
      write_address_data_log_force[3890] <= 6'h00;
      write_address_data_log_force[3891] <= 6'h00;
      write_address_data_log_force[3892] <= 6'h00;
      write_address_data_log_force[3893] <= 6'h00;
      write_address_data_log_force[3894] <= 6'h00;
      write_address_data_log_force[3895] <= 6'h00;
      write_address_data_log_force[3896] <= 6'h00;
      write_address_data_log_force[3897] <= 6'h00;
      write_address_data_log_force[3898] <= 6'h00;
      write_address_data_log_force[3899] <= 6'h00;
      write_address_data_log_force[3900] <= 6'h00;
      write_address_data_log_force[3901] <= 6'h00;
      write_address_data_log_force[3902] <= 6'h00;
      write_address_data_log_force[3903] <= 6'h00;
      write_address_data_log_force[3904] <= 6'h00;
      write_address_data_log_force[3905] <= 6'h00;
      write_address_data_log_force[3906] <= 6'h00;
      write_address_data_log_force[3907] <= 6'h00;
      write_address_data_log_force[3908] <= 6'h00;
      write_address_data_log_force[3909] <= 6'h00;
      write_address_data_log_force[3910] <= 6'h00;
      write_address_data_log_force[3911] <= 6'h00;
      write_address_data_log_force[3912] <= 6'h00;
      write_address_data_log_force[3913] <= 6'h00;
      write_address_data_log_force[3914] <= 6'h00;
      write_address_data_log_force[3915] <= 6'h00;
      write_address_data_log_force[3916] <= 6'h00;
      write_address_data_log_force[3917] <= 6'h00;
      write_address_data_log_force[3918] <= 6'h00;
      write_address_data_log_force[3919] <= 6'h00;
      write_address_data_log_force[3920] <= 6'h00;
      write_address_data_log_force[3921] <= 6'h00;
      write_address_data_log_force[3922] <= 6'h00;
      write_address_data_log_force[3923] <= 6'h00;
      write_address_data_log_force[3924] <= 6'h00;
      write_address_data_log_force[3925] <= 6'h00;
      write_address_data_log_force[3926] <= 6'h00;
      write_address_data_log_force[3927] <= 6'h00;
      write_address_data_log_force[3928] <= 6'h00;
      write_address_data_log_force[3929] <= 6'h00;
      write_address_data_log_force[3930] <= 6'h00;
      write_address_data_log_force[3931] <= 6'h00;
      write_address_data_log_force[3932] <= 6'h00;
      write_address_data_log_force[3933] <= 6'h00;
      write_address_data_log_force[3934] <= 6'h00;
      write_address_data_log_force[3935] <= 6'h00;
      write_address_data_log_force[3936] <= 6'h00;
      write_address_data_log_force[3937] <= 6'h00;
      write_address_data_log_force[3938] <= 6'h00;
      write_address_data_log_force[3939] <= 6'h00;
      write_address_data_log_force[3940] <= 6'h00;
      write_address_data_log_force[3941] <= 6'h00;
      write_address_data_log_force[3942] <= 6'h00;
      write_address_data_log_force[3943] <= 6'h00;
      write_address_data_log_force[3944] <= 6'h00;
      write_address_data_log_force[3945] <= 6'h00;
      write_address_data_log_force[3946] <= 6'h00;
      write_address_data_log_force[3947] <= 6'h00;
      write_address_data_log_force[3948] <= 6'h00;
      write_address_data_log_force[3949] <= 6'h00;
      write_address_data_log_force[3950] <= 6'h00;
      write_address_data_log_force[3951] <= 6'h00;
      write_address_data_log_force[3952] <= 6'h00;
      write_address_data_log_force[3953] <= 6'h00;
      write_address_data_log_force[3954] <= 6'h00;
      write_address_data_log_force[3955] <= 6'h00;
      write_address_data_log_force[3956] <= 6'h00;
      write_address_data_log_force[3957] <= 6'h00;
      write_address_data_log_force[3958] <= 6'h00;
      write_address_data_log_force[3959] <= 6'h00;
      write_address_data_log_force[3960] <= 6'h00;
      write_address_data_log_force[3961] <= 6'h00;
      write_address_data_log_force[3962] <= 6'h00;
      write_address_data_log_force[3963] <= 6'h00;
      write_address_data_log_force[3964] <= 6'h00;
      write_address_data_log_force[3965] <= 6'h00;
      write_address_data_log_force[3966] <= 6'h00;
      write_address_data_log_force[3967] <= 6'h00;
      write_address_data_log_force[3968] <= 6'h00;
      write_address_data_log_force[3969] <= 6'h00;
      write_address_data_log_force[3970] <= 6'h00;
      write_address_data_log_force[3971] <= 6'h00;
      write_address_data_log_force[3972] <= 6'h00;
      write_address_data_log_force[3973] <= 6'h00;
      write_address_data_log_force[3974] <= 6'h00;
      write_address_data_log_force[3975] <= 6'h00;
      write_address_data_log_force[3976] <= 6'h00;
      write_address_data_log_force[3977] <= 6'h00;
      write_address_data_log_force[3978] <= 6'h00;
      write_address_data_log_force[3979] <= 6'h00;
      write_address_data_log_force[3980] <= 6'h00;
      write_address_data_log_force[3981] <= 6'h00;
      write_address_data_log_force[3982] <= 6'h00;
      write_address_data_log_force[3983] <= 6'h00;
      write_address_data_log_force[3984] <= 6'h00;
      write_address_data_log_force[3985] <= 6'h00;
      write_address_data_log_force[3986] <= 6'h00;
      write_address_data_log_force[3987] <= 6'h00;
      write_address_data_log_force[3988] <= 6'h00;
      write_address_data_log_force[3989] <= 6'h00;
      write_address_data_log_force[3990] <= 6'h00;
      write_address_data_log_force[3991] <= 6'h00;
      write_address_data_log_force[3992] <= 6'h00;
      write_address_data_log_force[3993] <= 6'h00;
      write_address_data_log_force[3994] <= 6'h00;
      write_address_data_log_force[3995] <= 6'h00;
      write_address_data_log_force[3996] <= 6'h00;
      write_address_data_log_force[3997] <= 6'h00;
      write_address_data_log_force[3998] <= 6'h00;
      write_address_data_log_force[3999] <= 6'h00;
      write_address_data_log_force[4000] <= 6'h00;
      write_address_data_log_force[4001] <= 6'h00;
      write_address_data_log_force[4002] <= 6'h00;
      write_address_data_log_force[4003] <= 6'h00;
      write_address_data_log_force[4004] <= 6'h00;
      write_address_data_log_force[4005] <= 6'h00;
      write_address_data_log_force[4006] <= 6'h00;
      write_address_data_log_force[4007] <= 6'h00;
      write_address_data_log_force[4008] <= 6'h00;
      write_address_data_log_force[4009] <= 6'h00;
      write_address_data_log_force[4010] <= 6'h00;
      write_address_data_log_force[4011] <= 6'h00;
      write_address_data_log_force[4012] <= 6'h00;
      write_address_data_log_force[4013] <= 6'h00;
      write_address_data_log_force[4014] <= 6'h00;
      write_address_data_log_force[4015] <= 6'h00;
      write_address_data_log_force[4016] <= 6'h00;
      write_address_data_log_force[4017] <= 6'h00;
      write_address_data_log_force[4018] <= 6'h00;
      write_address_data_log_force[4019] <= 6'h00;
      write_address_data_log_force[4020] <= 6'h00;
      write_address_data_log_force[4021] <= 6'h00;
      write_address_data_log_force[4022] <= 6'h00;
      write_address_data_log_force[4023] <= 6'h00;
      write_address_data_log_force[4024] <= 6'h00;
      write_address_data_log_force[4025] <= 6'h00;
      write_address_data_log_force[4026] <= 6'h00;
      write_address_data_log_force[4027] <= 6'h00;
      write_address_data_log_force[4028] <= 6'h00;
      write_address_data_log_force[4029] <= 6'h00;
      write_address_data_log_force[4030] <= 6'h00;
      write_address_data_log_force[4031] <= 6'h00;
      write_address_data_log_force[4032] <= 6'h00;
      write_address_data_log_force[4033] <= 6'h00;
      write_address_data_log_force[4034] <= 6'h00;
      write_address_data_log_force[4035] <= 6'h00;
      write_address_data_log_force[4036] <= 6'h00;
      write_address_data_log_force[4037] <= 6'h00;
      write_address_data_log_force[4038] <= 6'h00;
      write_address_data_log_force[4039] <= 6'h00;
      write_address_data_log_force[4040] <= 6'h00;
      write_address_data_log_force[4041] <= 6'h00;
      write_address_data_log_force[4042] <= 6'h00;
      write_address_data_log_force[4043] <= 6'h00;
      write_address_data_log_force[4044] <= 6'h00;
      write_address_data_log_force[4045] <= 6'h00;
      write_address_data_log_force[4046] <= 6'h00;
      write_address_data_log_force[4047] <= 6'h00;
      write_address_data_log_force[4048] <= 6'h00;
      write_address_data_log_force[4049] <= 6'h00;
      write_address_data_log_force[4050] <= 6'h00;
      write_address_data_log_force[4051] <= 6'h00;
      write_address_data_log_force[4052] <= 6'h00;
      write_address_data_log_force[4053] <= 6'h00;
      write_address_data_log_force[4054] <= 6'h00;
      write_address_data_log_force[4055] <= 6'h00;
      write_address_data_log_force[4056] <= 6'h00;
      write_address_data_log_force[4057] <= 6'h00;
      write_address_data_log_force[4058] <= 6'h00;
      write_address_data_log_force[4059] <= 6'h00;
      write_address_data_log_force[4060] <= 6'h00;
      write_address_data_log_force[4061] <= 6'h00;
      write_address_data_log_force[4062] <= 6'h00;
      write_address_data_log_force[4063] <= 6'h00;
      write_address_data_log_force[4064] <= 6'h00;
      write_address_data_log_force[4065] <= 6'h00;
      write_address_data_log_force[4066] <= 6'h00;
      write_address_data_log_force[4067] <= 6'h00;
      write_address_data_log_force[4068] <= 6'h00;
      write_address_data_log_force[4069] <= 6'h00;
      write_address_data_log_force[4070] <= 6'h00;
      write_address_data_log_force[4071] <= 6'h00;
      write_address_data_log_force[4072] <= 6'h00;
      write_address_data_log_force[4073] <= 6'h00;
      write_address_data_log_force[4074] <= 6'h00;
      write_address_data_log_force[4075] <= 6'h00;
      write_address_data_log_force[4076] <= 6'h00;
      write_address_data_log_force[4077] <= 6'h00;
      write_address_data_log_force[4078] <= 6'h00;
      write_address_data_log_force[4079] <= 6'h00;
      write_address_data_log_force[4080] <= 6'h00;
      write_address_data_log_force[4081] <= 6'h00;
      write_address_data_log_force[4082] <= 6'h00;
      write_address_data_log_force[4083] <= 6'h00;
      write_address_data_log_force[4084] <= 6'h00;
      write_address_data_log_force[4085] <= 6'h00;
      write_address_data_log_force[4086] <= 6'h00;
      write_address_data_log_force[4087] <= 6'h00;
      write_address_data_log_force[4088] <= 6'h00;
      write_address_data_log_force[4089] <= 6'h00;
      write_address_data_log_force[4090] <= 6'h00;
      write_address_data_log_force[4091] <= 6'h00;
      write_address_data_log_force[4092] <= 6'h00;
      write_address_data_log_force[4093] <= 6'h00;
      write_address_data_log_force[4094] <= 6'h00;
      write_address_data_log_force[4095] <= 6'h00;
      write_address_data_log_force[4096] <= 6'h00;
      write_address_data_log_force[4097] <= 6'h00;
      write_address_data_log_force[4098] <= 6'h00;
      write_address_data_log_force[4099] <= 6'h00;
      write_address_data_log_force[4100] <= 6'h00;
      write_address_data_log_force[4101] <= 6'h00;
      write_address_data_log_force[4102] <= 6'h00;
      write_address_data_log_force[4103] <= 6'h00;
      write_address_data_log_force[4104] <= 6'h00;
      write_address_data_log_force[4105] <= 6'h00;
      write_address_data_log_force[4106] <= 6'h00;
      write_address_data_log_force[4107] <= 6'h00;
      write_address_data_log_force[4108] <= 6'h00;
      write_address_data_log_force[4109] <= 6'h00;
      write_address_data_log_force[4110] <= 6'h00;
      write_address_data_log_force[4111] <= 6'h00;
      write_address_data_log_force[4112] <= 6'h00;
      write_address_data_log_force[4113] <= 6'h00;
      write_address_data_log_force[4114] <= 6'h00;
      write_address_data_log_force[4115] <= 6'h00;
      write_address_data_log_force[4116] <= 6'h00;
      write_address_data_log_force[4117] <= 6'h00;
      write_address_data_log_force[4118] <= 6'h00;
      write_address_data_log_force[4119] <= 6'h00;
      write_address_data_log_force[4120] <= 6'h00;
      write_address_data_log_force[4121] <= 6'h00;
      write_address_data_log_force[4122] <= 6'h00;
      write_address_data_log_force[4123] <= 6'h00;
      write_address_data_log_force[4124] <= 6'h00;
      write_address_data_log_force[4125] <= 6'h00;
      write_address_data_log_force[4126] <= 6'h00;
      write_address_data_log_force[4127] <= 6'h00;
      write_address_data_log_force[4128] <= 6'h00;
      write_address_data_log_force[4129] <= 6'h00;
      write_address_data_log_force[4130] <= 6'h00;
      write_address_data_log_force[4131] <= 6'h00;
      write_address_data_log_force[4132] <= 6'h00;
      write_address_data_log_force[4133] <= 6'h00;
      write_address_data_log_force[4134] <= 6'h00;
      write_address_data_log_force[4135] <= 6'h00;
      write_address_data_log_force[4136] <= 6'h00;
      write_address_data_log_force[4137] <= 6'h00;
      write_address_data_log_force[4138] <= 6'h00;
      write_address_data_log_force[4139] <= 6'h00;
      write_address_data_log_force[4140] <= 6'h00;
      write_address_data_log_force[4141] <= 6'h00;
      write_address_data_log_force[4142] <= 6'h00;
      write_address_data_log_force[4143] <= 6'h00;
      write_address_data_log_force[4144] <= 6'h00;
      write_address_data_log_force[4145] <= 6'h00;
      write_address_data_log_force[4146] <= 6'h00;
      write_address_data_log_force[4147] <= 6'h00;
      write_address_data_log_force[4148] <= 6'h00;
      write_address_data_log_force[4149] <= 6'h00;
      write_address_data_log_force[4150] <= 6'h00;
      write_address_data_log_force[4151] <= 6'h00;
      write_address_data_log_force[4152] <= 6'h00;
      write_address_data_log_force[4153] <= 6'h00;
      write_address_data_log_force[4154] <= 6'h00;
      write_address_data_log_force[4155] <= 6'h00;
      write_address_data_log_force[4156] <= 6'h00;
      write_address_data_log_force[4157] <= 6'h00;
      write_address_data_log_force[4158] <= 6'h00;
      write_address_data_log_force[4159] <= 6'h00;
      write_address_data_log_force[4160] <= 6'h00;
      write_address_data_log_force[4161] <= 6'h00;
      write_address_data_log_force[4162] <= 6'h00;
      write_address_data_log_force[4163] <= 6'h00;
      write_address_data_log_force[4164] <= 6'h00;
      write_address_data_log_force[4165] <= 6'h00;
      write_address_data_log_force[4166] <= 6'h00;
      write_address_data_log_force[4167] <= 6'h00;
      write_address_data_log_force[4168] <= 6'h00;
      write_address_data_log_force[4169] <= 6'h00;
      write_address_data_log_force[4170] <= 6'h00;
      write_address_data_log_force[4171] <= 6'h00;
      write_address_data_log_force[4172] <= 6'h00;
      write_address_data_log_force[4173] <= 6'h00;
      write_address_data_log_force[4174] <= 6'h00;
      write_address_data_log_force[4175] <= 6'h00;
      write_address_data_log_force[4176] <= 6'h00;
      write_address_data_log_force[4177] <= 6'h00;
      write_address_data_log_force[4178] <= 6'h00;
      write_address_data_log_force[4179] <= 6'h00;
      write_address_data_log_force[4180] <= 6'h00;
      write_address_data_log_force[4181] <= 6'h00;
      write_address_data_log_force[4182] <= 6'h00;
      write_address_data_log_force[4183] <= 6'h00;
      write_address_data_log_force[4184] <= 6'h00;
      write_address_data_log_force[4185] <= 6'h00;
      write_address_data_log_force[4186] <= 6'h00;
      write_address_data_log_force[4187] <= 6'h00;
      write_address_data_log_force[4188] <= 6'h00;
      write_address_data_log_force[4189] <= 6'h00;
      write_address_data_log_force[4190] <= 6'h00;
      write_address_data_log_force[4191] <= 6'h00;
      write_address_data_log_force[4192] <= 6'h00;
      write_address_data_log_force[4193] <= 6'h00;
      write_address_data_log_force[4194] <= 6'h00;
      write_address_data_log_force[4195] <= 6'h00;
      write_address_data_log_force[4196] <= 6'h00;
      write_address_data_log_force[4197] <= 6'h00;
      write_address_data_log_force[4198] <= 6'h00;
      write_address_data_log_force[4199] <= 6'h00;
      write_address_data_log_force[4200] <= 6'h00;
      write_address_data_log_force[4201] <= 6'h00;
      write_address_data_log_force[4202] <= 6'h00;
      write_address_data_log_force[4203] <= 6'h00;
      write_address_data_log_force[4204] <= 6'h00;
      write_address_data_log_force[4205] <= 6'h00;
      write_address_data_log_force[4206] <= 6'h00;
      write_address_data_log_force[4207] <= 6'h00;
      write_address_data_log_force[4208] <= 6'h00;
      write_address_data_log_force[4209] <= 6'h00;
      write_address_data_log_force[4210] <= 6'h00;
      write_address_data_log_force[4211] <= 6'h00;
      write_address_data_log_force[4212] <= 6'h00;
      write_address_data_log_force[4213] <= 6'h00;
      write_address_data_log_force[4214] <= 6'h00;
      write_address_data_log_force[4215] <= 6'h00;
      write_address_data_log_force[4216] <= 6'h00;
      write_address_data_log_force[4217] <= 6'h00;
      write_address_data_log_force[4218] <= 6'h00;
      write_address_data_log_force[4219] <= 6'h00;
      write_address_data_log_force[4220] <= 6'h00;
      write_address_data_log_force[4221] <= 6'h00;
      write_address_data_log_force[4222] <= 6'h00;
      write_address_data_log_force[4223] <= 6'h00;
      write_address_data_log_force[4224] <= 6'h00;
      write_address_data_log_force[4225] <= 6'h00;
      write_address_data_log_force[4226] <= 6'h00;
      write_address_data_log_force[4227] <= 6'h00;
      write_address_data_log_force[4228] <= 6'h00;
      write_address_data_log_force[4229] <= 6'h00;
      write_address_data_log_force[4230] <= 6'h00;
      write_address_data_log_force[4231] <= 6'h00;
      write_address_data_log_force[4232] <= 6'h00;
      write_address_data_log_force[4233] <= 6'h00;
      write_address_data_log_force[4234] <= 6'h00;
      write_address_data_log_force[4235] <= 6'h00;
      write_address_data_log_force[4236] <= 6'h00;
      write_address_data_log_force[4237] <= 6'h00;
      write_address_data_log_force[4238] <= 6'h00;
      write_address_data_log_force[4239] <= 6'h00;
      write_address_data_log_force[4240] <= 6'h00;
      write_address_data_log_force[4241] <= 6'h00;
      write_address_data_log_force[4242] <= 6'h00;
      write_address_data_log_force[4243] <= 6'h00;
      write_address_data_log_force[4244] <= 6'h00;
      write_address_data_log_force[4245] <= 6'h00;
      write_address_data_log_force[4246] <= 6'h00;
      write_address_data_log_force[4247] <= 6'h00;
      write_address_data_log_force[4248] <= 6'h00;
      write_address_data_log_force[4249] <= 6'h00;
      write_address_data_log_force[4250] <= 6'h00;
      write_address_data_log_force[4251] <= 6'h00;
      write_address_data_log_force[4252] <= 6'h00;
      write_address_data_log_force[4253] <= 6'h00;
      write_address_data_log_force[4254] <= 6'h00;
      write_address_data_log_force[4255] <= 6'h00;
      write_address_data_log_force[4256] <= 6'h00;
      write_address_data_log_force[4257] <= 6'h00;
      write_address_data_log_force[4258] <= 6'h00;
      write_address_data_log_force[4259] <= 6'h00;
      write_address_data_log_force[4260] <= 6'h00;
      write_address_data_log_force[4261] <= 6'h00;
      write_address_data_log_force[4262] <= 6'h00;
      write_address_data_log_force[4263] <= 6'h00;
      write_address_data_log_force[4264] <= 6'h00;
      write_address_data_log_force[4265] <= 6'h00;
      write_address_data_log_force[4266] <= 6'h00;
      write_address_data_log_force[4267] <= 6'h00;
      write_address_data_log_force[4268] <= 6'h00;
      write_address_data_log_force[4269] <= 6'h00;
      write_address_data_log_force[4270] <= 6'h00;
      write_address_data_log_force[4271] <= 6'h00;
      write_address_data_log_force[4272] <= 6'h00;
      write_address_data_log_force[4273] <= 6'h00;
      write_address_data_log_force[4274] <= 6'h00;
      write_address_data_log_force[4275] <= 6'h00;
      write_address_data_log_force[4276] <= 6'h00;
      write_address_data_log_force[4277] <= 6'h00;
      write_address_data_log_force[4278] <= 6'h00;
      write_address_data_log_force[4279] <= 6'h00;
      write_address_data_log_force[4280] <= 6'h00;
      write_address_data_log_force[4281] <= 6'h00;
      write_address_data_log_force[4282] <= 6'h00;
      write_address_data_log_force[4283] <= 6'h00;
      write_address_data_log_force[4284] <= 6'h00;
      write_address_data_log_force[4285] <= 6'h00;
      write_address_data_log_force[4286] <= 6'h00;
      write_address_data_log_force[4287] <= 6'h00;
      write_address_data_log_force[4288] <= 6'h00;
      write_address_data_log_force[4289] <= 6'h00;
      write_address_data_log_force[4290] <= 6'h00;
      write_address_data_log_force[4291] <= 6'h00;
      write_address_data_log_force[4292] <= 6'h00;
      write_address_data_log_force[4293] <= 6'h00;
      write_address_data_log_force[4294] <= 6'h00;
      write_address_data_log_force[4295] <= 6'h00;
      write_address_data_log_force[4296] <= 6'h00;
      write_address_data_log_force[4297] <= 6'h00;
      write_address_data_log_force[4298] <= 6'h00;
      write_address_data_log_force[4299] <= 6'h00;
      write_address_data_log_force[4300] <= 6'h00;
      write_address_data_log_force[4301] <= 6'h00;
      write_address_data_log_force[4302] <= 6'h00;
      write_address_data_log_force[4303] <= 6'h00;
      write_address_data_log_force[4304] <= 6'h00;
      write_address_data_log_force[4305] <= 6'h00;
      write_address_data_log_force[4306] <= 6'h00;
      write_address_data_log_force[4307] <= 6'h00;
      write_address_data_log_force[4308] <= 6'h00;
      write_address_data_log_force[4309] <= 6'h00;
      write_address_data_log_force[4310] <= 6'h00;
      write_address_data_log_force[4311] <= 6'h00;
      write_address_data_log_force[4312] <= 6'h00;
      write_address_data_log_force[4313] <= 6'h00;
      write_address_data_log_force[4314] <= 6'h00;
      write_address_data_log_force[4315] <= 6'h00;
      write_address_data_log_force[4316] <= 6'h00;
      write_address_data_log_force[4317] <= 6'h00;
      write_address_data_log_force[4318] <= 6'h00;
      write_address_data_log_force[4319] <= 6'h00;
      write_address_data_log_force[4320] <= 6'h00;
      write_address_data_log_force[4321] <= 6'h00;
      write_address_data_log_force[4322] <= 6'h00;
      write_address_data_log_force[4323] <= 6'h00;
      write_address_data_log_force[4324] <= 6'h00;
      write_address_data_log_force[4325] <= 6'h00;
      write_address_data_log_force[4326] <= 6'h00;
      write_address_data_log_force[4327] <= 6'h00;
      write_address_data_log_force[4328] <= 6'h00;
      write_address_data_log_force[4329] <= 6'h00;
      write_address_data_log_force[4330] <= 6'h00;
      write_address_data_log_force[4331] <= 6'h00;
      write_address_data_log_force[4332] <= 6'h00;
      write_address_data_log_force[4333] <= 6'h00;
      write_address_data_log_force[4334] <= 6'h00;
      write_address_data_log_force[4335] <= 6'h00;
      write_address_data_log_force[4336] <= 6'h00;
      write_address_data_log_force[4337] <= 6'h00;
      write_address_data_log_force[4338] <= 6'h00;
      write_address_data_log_force[4339] <= 6'h00;
      write_address_data_log_force[4340] <= 6'h00;
      write_address_data_log_force[4341] <= 6'h00;
      write_address_data_log_force[4342] <= 6'h00;
      write_address_data_log_force[4343] <= 6'h00;
      write_address_data_log_force[4344] <= 6'h00;
      write_address_data_log_force[4345] <= 6'h00;
      write_address_data_log_force[4346] <= 6'h00;
      write_address_data_log_force[4347] <= 6'h00;
      write_address_data_log_force[4348] <= 6'h00;
      write_address_data_log_force[4349] <= 6'h00;
      write_address_data_log_force[4350] <= 6'h00;
      write_address_data_log_force[4351] <= 6'h00;
      write_address_data_log_force[4352] <= 6'h00;
      write_address_data_log_force[4353] <= 6'h00;
      write_address_data_log_force[4354] <= 6'h00;
      write_address_data_log_force[4355] <= 6'h00;
      write_address_data_log_force[4356] <= 6'h00;
      write_address_data_log_force[4357] <= 6'h00;
      write_address_data_log_force[4358] <= 6'h00;
      write_address_data_log_force[4359] <= 6'h00;
      write_address_data_log_force[4360] <= 6'h00;
      write_address_data_log_force[4361] <= 6'h00;
      write_address_data_log_force[4362] <= 6'h00;
      write_address_data_log_force[4363] <= 6'h00;
      write_address_data_log_force[4364] <= 6'h00;
      write_address_data_log_force[4365] <= 6'h00;
      write_address_data_log_force[4366] <= 6'h00;
      write_address_data_log_force[4367] <= 6'h00;
      write_address_data_log_force[4368] <= 6'h00;
      write_address_data_log_force[4369] <= 6'h00;
      write_address_data_log_force[4370] <= 6'h00;
      write_address_data_log_force[4371] <= 6'h00;
      write_address_data_log_force[4372] <= 6'h00;
      write_address_data_log_force[4373] <= 6'h00;
      write_address_data_log_force[4374] <= 6'h00;
      write_address_data_log_force[4375] <= 6'h00;
      write_address_data_log_force[4376] <= 6'h00;
      write_address_data_log_force[4377] <= 6'h00;
      write_address_data_log_force[4378] <= 6'h00;
      write_address_data_log_force[4379] <= 6'h00;
      write_address_data_log_force[4380] <= 6'h00;
      write_address_data_log_force[4381] <= 6'h00;
      write_address_data_log_force[4382] <= 6'h00;
      write_address_data_log_force[4383] <= 6'h00;
      write_address_data_log_force[4384] <= 6'h00;
      write_address_data_log_force[4385] <= 6'h00;
      write_address_data_log_force[4386] <= 6'h00;
      write_address_data_log_force[4387] <= 6'h00;
      write_address_data_log_force[4388] <= 6'h00;
      write_address_data_log_force[4389] <= 6'h00;
      write_address_data_log_force[4390] <= 6'h00;
      write_address_data_log_force[4391] <= 6'h00;
      write_address_data_log_force[4392] <= 6'h00;
      write_address_data_log_force[4393] <= 6'h00;
      write_address_data_log_force[4394] <= 6'h00;
      write_address_data_log_force[4395] <= 6'h00;
      write_address_data_log_force[4396] <= 6'h00;
      write_address_data_log_force[4397] <= 6'h00;
      write_address_data_log_force[4398] <= 6'h00;
      write_address_data_log_force[4399] <= 6'h00;
      write_address_data_log_force[4400] <= 6'h00;
      write_address_data_log_force[4401] <= 6'h00;
      write_address_data_log_force[4402] <= 6'h00;
      write_address_data_log_force[4403] <= 6'h00;
      write_address_data_log_force[4404] <= 6'h00;
      write_address_data_log_force[4405] <= 6'h00;
      write_address_data_log_force[4406] <= 6'h00;
      write_address_data_log_force[4407] <= 6'h00;
      write_address_data_log_force[4408] <= 6'h00;
      write_address_data_log_force[4409] <= 6'h00;
      write_address_data_log_force[4410] <= 6'h00;
      write_address_data_log_force[4411] <= 6'h00;
      write_address_data_log_force[4412] <= 6'h00;
      write_address_data_log_force[4413] <= 6'h00;
      write_address_data_log_force[4414] <= 6'h00;
      write_address_data_log_force[4415] <= 6'h00;
      write_address_data_log_force[4416] <= 6'h00;
      write_address_data_log_force[4417] <= 6'h00;
      write_address_data_log_force[4418] <= 6'h00;
      write_address_data_log_force[4419] <= 6'h00;
      write_address_data_log_force[4420] <= 6'h00;
      write_address_data_log_force[4421] <= 6'h00;
      write_address_data_log_force[4422] <= 6'h00;
      write_address_data_log_force[4423] <= 6'h00;
      write_address_data_log_force[4424] <= 6'h00;
      write_address_data_log_force[4425] <= 6'h00;
      write_address_data_log_force[4426] <= 6'h00;
      write_address_data_log_force[4427] <= 6'h00;
      write_address_data_log_force[4428] <= 6'h00;
      write_address_data_log_force[4429] <= 6'h00;
      write_address_data_log_force[4430] <= 6'h00;
      write_address_data_log_force[4431] <= 6'h00;
      write_address_data_log_force[4432] <= 6'h00;
      write_address_data_log_force[4433] <= 6'h00;
      write_address_data_log_force[4434] <= 6'h00;
      write_address_data_log_force[4435] <= 6'h00;
      write_address_data_log_force[4436] <= 6'h00;
      write_address_data_log_force[4437] <= 6'h00;
      write_address_data_log_force[4438] <= 6'h00;
      write_address_data_log_force[4439] <= 6'h00;
      write_address_data_log_force[4440] <= 6'h00;
      write_address_data_log_force[4441] <= 6'h00;
      write_address_data_log_force[4442] <= 6'h00;
      write_address_data_log_force[4443] <= 6'h00;
      write_address_data_log_force[4444] <= 6'h00;
      write_address_data_log_force[4445] <= 6'h00;
      write_address_data_log_force[4446] <= 6'h00;
      write_address_data_log_force[4447] <= 6'h00;
      write_address_data_log_force[4448] <= 6'h00;
      write_address_data_log_force[4449] <= 6'h00;
      write_address_data_log_force[4450] <= 6'h00;
      write_address_data_log_force[4451] <= 6'h00;
      write_address_data_log_force[4452] <= 6'h00;
      write_address_data_log_force[4453] <= 6'h00;
      write_address_data_log_force[4454] <= 6'h00;
      write_address_data_log_force[4455] <= 6'h00;
      write_address_data_log_force[4456] <= 6'h00;
      write_address_data_log_force[4457] <= 6'h00;
      write_address_data_log_force[4458] <= 6'h00;
      write_address_data_log_force[4459] <= 6'h00;
      write_address_data_log_force[4460] <= 6'h00;
      write_address_data_log_force[4461] <= 6'h00;
      write_address_data_log_force[4462] <= 6'h00;
      write_address_data_log_force[4463] <= 6'h00;
      write_address_data_log_force[4464] <= 6'h00;
      write_address_data_log_force[4465] <= 6'h00;
      write_address_data_log_force[4466] <= 6'h00;
      write_address_data_log_force[4467] <= 6'h00;
      write_address_data_log_force[4468] <= 6'h00;
      write_address_data_log_force[4469] <= 6'h00;
      write_address_data_log_force[4470] <= 6'h00;
      write_address_data_log_force[4471] <= 6'h00;
      write_address_data_log_force[4472] <= 6'h00;
      write_address_data_log_force[4473] <= 6'h00;
      write_address_data_log_force[4474] <= 6'h00;
      write_address_data_log_force[4475] <= 6'h00;
      write_address_data_log_force[4476] <= 6'h00;
      write_address_data_log_force[4477] <= 6'h00;
      write_address_data_log_force[4478] <= 6'h00;
      write_address_data_log_force[4479] <= 6'h00;
      write_address_data_log_force[4480] <= 6'h00;
      write_address_data_log_force[4481] <= 6'h00;
      write_address_data_log_force[4482] <= 6'h00;
      write_address_data_log_force[4483] <= 6'h00;
      write_address_data_log_force[4484] <= 6'h00;
      write_address_data_log_force[4485] <= 6'h00;
      write_address_data_log_force[4486] <= 6'h00;
      write_address_data_log_force[4487] <= 6'h00;
      write_address_data_log_force[4488] <= 6'h00;
      write_address_data_log_force[4489] <= 6'h00;
      write_address_data_log_force[4490] <= 6'h00;
      write_address_data_log_force[4491] <= 6'h00;
      write_address_data_log_force[4492] <= 6'h00;
      write_address_data_log_force[4493] <= 6'h00;
      write_address_data_log_force[4494] <= 6'h00;
      write_address_data_log_force[4495] <= 6'h00;
      write_address_data_log_force[4496] <= 6'h00;
      write_address_data_log_force[4497] <= 6'h00;
      write_address_data_log_force[4498] <= 6'h00;
      write_address_data_log_force[4499] <= 6'h00;
      write_address_data_log_force[4500] <= 6'h00;
      write_address_data_log_force[4501] <= 6'h00;
      write_address_data_log_force[4502] <= 6'h00;
      write_address_data_log_force[4503] <= 6'h00;
      write_address_data_log_force[4504] <= 6'h00;
      write_address_data_log_force[4505] <= 6'h00;
      write_address_data_log_force[4506] <= 6'h00;
      write_address_data_log_force[4507] <= 6'h00;
      write_address_data_log_force[4508] <= 6'h00;
      write_address_data_log_force[4509] <= 6'h00;
      write_address_data_log_force[4510] <= 6'h00;
      write_address_data_log_force[4511] <= 6'h00;
      write_address_data_log_force[4512] <= 6'h00;
      write_address_data_log_force[4513] <= 6'h00;
      write_address_data_log_force[4514] <= 6'h00;
      write_address_data_log_force[4515] <= 6'h00;
      write_address_data_log_force[4516] <= 6'h00;
      write_address_data_log_force[4517] <= 6'h00;
      write_address_data_log_force[4518] <= 6'h00;
      write_address_data_log_force[4519] <= 6'h00;
      write_address_data_log_force[4520] <= 6'h00;
      write_address_data_log_force[4521] <= 6'h00;
      write_address_data_log_force[4522] <= 6'h00;
      write_address_data_log_force[4523] <= 6'h00;
      write_address_data_log_force[4524] <= 6'h00;
      write_address_data_log_force[4525] <= 6'h00;
      write_address_data_log_force[4526] <= 6'h00;
      write_address_data_log_force[4527] <= 6'h00;
      write_address_data_log_force[4528] <= 6'h00;
      write_address_data_log_force[4529] <= 6'h00;
      write_address_data_log_force[4530] <= 6'h00;
      write_address_data_log_force[4531] <= 6'h00;
      write_address_data_log_force[4532] <= 6'h00;
      write_address_data_log_force[4533] <= 6'h00;
      write_address_data_log_force[4534] <= 6'h00;
      write_address_data_log_force[4535] <= 6'h00;
      write_address_data_log_force[4536] <= 6'h00;
      write_address_data_log_force[4537] <= 6'h00;
      write_address_data_log_force[4538] <= 6'h00;
      write_address_data_log_force[4539] <= 6'h00;
      write_address_data_log_force[4540] <= 6'h00;
      write_address_data_log_force[4541] <= 6'h00;
      write_address_data_log_force[4542] <= 6'h00;
      write_address_data_log_force[4543] <= 6'h00;
      write_address_data_log_force[4544] <= 6'h00;
      write_address_data_log_force[4545] <= 6'h00;
      write_address_data_log_force[4546] <= 6'h00;
      write_address_data_log_force[4547] <= 6'h00;
      write_address_data_log_force[4548] <= 6'h00;
      write_address_data_log_force[4549] <= 6'h00;
      write_address_data_log_force[4550] <= 6'h00;
      write_address_data_log_force[4551] <= 6'h00;
      write_address_data_log_force[4552] <= 6'h00;
      write_address_data_log_force[4553] <= 6'h00;
      write_address_data_log_force[4554] <= 6'h00;
      write_address_data_log_force[4555] <= 6'h00;
      write_address_data_log_force[4556] <= 6'h00;
      write_address_data_log_force[4557] <= 6'h00;
      write_address_data_log_force[4558] <= 6'h00;
      write_address_data_log_force[4559] <= 6'h00;
      write_address_data_log_force[4560] <= 6'h00;
      write_address_data_log_force[4561] <= 6'h00;
      write_address_data_log_force[4562] <= 6'h00;
      write_address_data_log_force[4563] <= 6'h00;
      write_address_data_log_force[4564] <= 6'h00;
      write_address_data_log_force[4565] <= 6'h00;
      write_address_data_log_force[4566] <= 6'h00;
      write_address_data_log_force[4567] <= 6'h00;
      write_address_data_log_force[4568] <= 6'h00;
      write_address_data_log_force[4569] <= 6'h00;
      write_address_data_log_force[4570] <= 6'h00;
      write_address_data_log_force[4571] <= 6'h00;
      write_address_data_log_force[4572] <= 6'h00;
      write_address_data_log_force[4573] <= 6'h00;
      write_address_data_log_force[4574] <= 6'h00;
      write_address_data_log_force[4575] <= 6'h00;
      write_address_data_log_force[4576] <= 6'h00;
      write_address_data_log_force[4577] <= 6'h00;
      write_address_data_log_force[4578] <= 6'h00;
      write_address_data_log_force[4579] <= 6'h00;
      write_address_data_log_force[4580] <= 6'h00;
      write_address_data_log_force[4581] <= 6'h00;
      write_address_data_log_force[4582] <= 6'h00;
      write_address_data_log_force[4583] <= 6'h00;
      write_address_data_log_force[4584] <= 6'h00;
      write_address_data_log_force[4585] <= 6'h00;
      write_address_data_log_force[4586] <= 6'h00;
      write_address_data_log_force[4587] <= 6'h00;
      write_address_data_log_force[4588] <= 6'h00;
      write_address_data_log_force[4589] <= 6'h00;
      write_address_data_log_force[4590] <= 6'h00;
      write_address_data_log_force[4591] <= 6'h00;
      write_address_data_log_force[4592] <= 6'h00;
      write_address_data_log_force[4593] <= 6'h00;
      write_address_data_log_force[4594] <= 6'h00;
      write_address_data_log_force[4595] <= 6'h00;
      write_address_data_log_force[4596] <= 6'h00;
      write_address_data_log_force[4597] <= 6'h00;
      write_address_data_log_force[4598] <= 6'h00;
      write_address_data_log_force[4599] <= 6'h00;
      write_address_data_log_force[4600] <= 6'h00;
      write_address_data_log_force[4601] <= 6'h00;
      write_address_data_log_force[4602] <= 6'h00;
      write_address_data_log_force[4603] <= 6'h00;
      write_address_data_log_force[4604] <= 6'h00;
      write_address_data_log_force[4605] <= 6'h00;
      write_address_data_log_force[4606] <= 6'h00;
      write_address_data_log_force[4607] <= 6'h00;
      write_address_data_log_force[4608] <= 6'h00;
      write_address_data_log_force[4609] <= 6'h00;
      write_address_data_log_force[4610] <= 6'h00;
      write_address_data_log_force[4611] <= 6'h00;
      write_address_data_log_force[4612] <= 6'h00;
      write_address_data_log_force[4613] <= 6'h00;
      write_address_data_log_force[4614] <= 6'h00;
      write_address_data_log_force[4615] <= 6'h00;
      write_address_data_log_force[4616] <= 6'h00;
      write_address_data_log_force[4617] <= 6'h00;
      write_address_data_log_force[4618] <= 6'h00;
      write_address_data_log_force[4619] <= 6'h00;
      write_address_data_log_force[4620] <= 6'h00;
      write_address_data_log_force[4621] <= 6'h00;
      write_address_data_log_force[4622] <= 6'h00;
      write_address_data_log_force[4623] <= 6'h00;
      write_address_data_log_force[4624] <= 6'h00;
      write_address_data_log_force[4625] <= 6'h00;
      write_address_data_log_force[4626] <= 6'h00;
      write_address_data_log_force[4627] <= 6'h00;
      write_address_data_log_force[4628] <= 6'h00;
      write_address_data_log_force[4629] <= 6'h00;
      write_address_data_log_force[4630] <= 6'h00;
      write_address_data_log_force[4631] <= 6'h00;
      write_address_data_log_force[4632] <= 6'h00;
      write_address_data_log_force[4633] <= 6'h00;
      write_address_data_log_force[4634] <= 6'h00;
      write_address_data_log_force[4635] <= 6'h00;
      write_address_data_log_force[4636] <= 6'h00;
      write_address_data_log_force[4637] <= 6'h00;
      write_address_data_log_force[4638] <= 6'h00;
      write_address_data_log_force[4639] <= 6'h00;
      write_address_data_log_force[4640] <= 6'h00;
      write_address_data_log_force[4641] <= 6'h00;
      write_address_data_log_force[4642] <= 6'h00;
      write_address_data_log_force[4643] <= 6'h00;
      write_address_data_log_force[4644] <= 6'h00;
      write_address_data_log_force[4645] <= 6'h00;
      write_address_data_log_force[4646] <= 6'h00;
      write_address_data_log_force[4647] <= 6'h00;
      write_address_data_log_force[4648] <= 6'h00;
      write_address_data_log_force[4649] <= 6'h00;
      write_address_data_log_force[4650] <= 6'h00;
      write_address_data_log_force[4651] <= 6'h00;
      write_address_data_log_force[4652] <= 6'h00;
      write_address_data_log_force[4653] <= 6'h00;
      write_address_data_log_force[4654] <= 6'h00;
      write_address_data_log_force[4655] <= 6'h00;
      write_address_data_log_force[4656] <= 6'h00;
      write_address_data_log_force[4657] <= 6'h00;
      write_address_data_log_force[4658] <= 6'h00;
      write_address_data_log_force[4659] <= 6'h00;
      write_address_data_log_force[4660] <= 6'h00;
      write_address_data_log_force[4661] <= 6'h00;
      write_address_data_log_force[4662] <= 6'h00;
      write_address_data_log_force[4663] <= 6'h00;
      write_address_data_log_force[4664] <= 6'h00;
      write_address_data_log_force[4665] <= 6'h00;
      write_address_data_log_force[4666] <= 6'h00;
      write_address_data_log_force[4667] <= 6'h00;
      write_address_data_log_force[4668] <= 6'h00;
      write_address_data_log_force[4669] <= 6'h00;
      write_address_data_log_force[4670] <= 6'h00;
      write_address_data_log_force[4671] <= 6'h00;
      write_address_data_log_force[4672] <= 6'h00;
      write_address_data_log_force[4673] <= 6'h00;
      write_address_data_log_force[4674] <= 6'h00;
      write_address_data_log_force[4675] <= 6'h00;
      write_address_data_log_force[4676] <= 6'h00;
      write_address_data_log_force[4677] <= 6'h00;
      write_address_data_log_force[4678] <= 6'h00;
      write_address_data_log_force[4679] <= 6'h00;
      write_address_data_log_force[4680] <= 6'h00;
      write_address_data_log_force[4681] <= 6'h00;
      write_address_data_log_force[4682] <= 6'h00;
      write_address_data_log_force[4683] <= 6'h00;
      write_address_data_log_force[4684] <= 6'h00;
      write_address_data_log_force[4685] <= 6'h00;
      write_address_data_log_force[4686] <= 6'h00;
      write_address_data_log_force[4687] <= 6'h00;
      write_address_data_log_force[4688] <= 6'h00;
      write_address_data_log_force[4689] <= 6'h00;
      write_address_data_log_force[4690] <= 6'h00;
      write_address_data_log_force[4691] <= 6'h00;
      write_address_data_log_force[4692] <= 6'h00;
      write_address_data_log_force[4693] <= 6'h00;
      write_address_data_log_force[4694] <= 6'h00;
      write_address_data_log_force[4695] <= 6'h00;
      write_address_data_log_force[4696] <= 6'h00;
      write_address_data_log_force[4697] <= 6'h00;
      write_address_data_log_force[4698] <= 6'h00;
      write_address_data_log_force[4699] <= 6'h00;
      write_address_data_log_force[4700] <= 6'h00;
      write_address_data_log_force[4701] <= 6'h00;
      write_address_data_log_force[4702] <= 6'h00;
      write_address_data_log_force[4703] <= 6'h00;
      write_address_data_log_force[4704] <= 6'h00;
      write_address_data_log_force[4705] <= 6'h00;
      write_address_data_log_force[4706] <= 6'h00;
      write_address_data_log_force[4707] <= 6'h00;
      write_address_data_log_force[4708] <= 6'h00;
      write_address_data_log_force[4709] <= 6'h00;
      write_address_data_log_force[4710] <= 6'h00;
      write_address_data_log_force[4711] <= 6'h00;
      write_address_data_log_force[4712] <= 6'h00;
      write_address_data_log_force[4713] <= 6'h00;
      write_address_data_log_force[4714] <= 6'h00;
      write_address_data_log_force[4715] <= 6'h00;
      write_address_data_log_force[4716] <= 6'h00;
      write_address_data_log_force[4717] <= 6'h00;
      write_address_data_log_force[4718] <= 6'h00;
      write_address_data_log_force[4719] <= 6'h00;
      write_address_data_log_force[4720] <= 6'h00;
      write_address_data_log_force[4721] <= 6'h00;
      write_address_data_log_force[4722] <= 6'h00;
      write_address_data_log_force[4723] <= 6'h00;
      write_address_data_log_force[4724] <= 6'h00;
      write_address_data_log_force[4725] <= 6'h00;
      write_address_data_log_force[4726] <= 6'h00;
      write_address_data_log_force[4727] <= 6'h00;
      write_address_data_log_force[4728] <= 6'h00;
      write_address_data_log_force[4729] <= 6'h00;
      write_address_data_log_force[4730] <= 6'h00;
      write_address_data_log_force[4731] <= 6'h00;
      write_address_data_log_force[4732] <= 6'h00;
      write_address_data_log_force[4733] <= 6'h00;
      write_address_data_log_force[4734] <= 6'h00;
      write_address_data_log_force[4735] <= 6'h00;
      write_address_data_log_force[4736] <= 6'h00;
      write_address_data_log_force[4737] <= 6'h00;
      write_address_data_log_force[4738] <= 6'h00;
      write_address_data_log_force[4739] <= 6'h00;
      write_address_data_log_force[4740] <= 6'h00;
      write_address_data_log_force[4741] <= 6'h00;
      write_address_data_log_force[4742] <= 6'h00;
      write_address_data_log_force[4743] <= 6'h00;
      write_address_data_log_force[4744] <= 6'h00;
      write_address_data_log_force[4745] <= 6'h00;
      write_address_data_log_force[4746] <= 6'h00;
      write_address_data_log_force[4747] <= 6'h00;
      write_address_data_log_force[4748] <= 6'h00;
      write_address_data_log_force[4749] <= 6'h00;
      write_address_data_log_force[4750] <= 6'h00;
      write_address_data_log_force[4751] <= 6'h00;
      write_address_data_log_force[4752] <= 6'h00;
      write_address_data_log_force[4753] <= 6'h00;
      write_address_data_log_force[4754] <= 6'h00;
      write_address_data_log_force[4755] <= 6'h00;
      write_address_data_log_force[4756] <= 6'h00;
      write_address_data_log_force[4757] <= 6'h00;
      write_address_data_log_force[4758] <= 6'h00;
      write_address_data_log_force[4759] <= 6'h00;
      write_address_data_log_force[4760] <= 6'h00;
      write_address_data_log_force[4761] <= 6'h00;
      write_address_data_log_force[4762] <= 6'h00;
      write_address_data_log_force[4763] <= 6'h00;
      write_address_data_log_force[4764] <= 6'h00;
      write_address_data_log_force[4765] <= 6'h00;
      write_address_data_log_force[4766] <= 6'h00;
      write_address_data_log_force[4767] <= 6'h00;
      write_address_data_log_force[4768] <= 6'h00;
      write_address_data_log_force[4769] <= 6'h00;
      write_address_data_log_force[4770] <= 6'h00;
      write_address_data_log_force[4771] <= 6'h00;
      write_address_data_log_force[4772] <= 6'h00;
      write_address_data_log_force[4773] <= 6'h00;
      write_address_data_log_force[4774] <= 6'h00;
      write_address_data_log_force[4775] <= 6'h00;
      write_address_data_log_force[4776] <= 6'h00;
      write_address_data_log_force[4777] <= 6'h00;
      write_address_data_log_force[4778] <= 6'h00;
      write_address_data_log_force[4779] <= 6'h00;
      write_address_data_log_force[4780] <= 6'h00;
      write_address_data_log_force[4781] <= 6'h00;
      write_address_data_log_force[4782] <= 6'h00;
      write_address_data_log_force[4783] <= 6'h00;
      write_address_data_log_force[4784] <= 6'h00;
      write_address_data_log_force[4785] <= 6'h00;
      write_address_data_log_force[4786] <= 6'h00;
      write_address_data_log_force[4787] <= 6'h00;
      write_address_data_log_force[4788] <= 6'h00;
      write_address_data_log_force[4789] <= 6'h00;
      write_address_data_log_force[4790] <= 6'h00;
      write_address_data_log_force[4791] <= 6'h00;
      write_address_data_log_force[4792] <= 6'h00;
      write_address_data_log_force[4793] <= 6'h00;
      write_address_data_log_force[4794] <= 6'h00;
      write_address_data_log_force[4795] <= 6'h00;
      write_address_data_log_force[4796] <= 6'h00;
      write_address_data_log_force[4797] <= 6'h00;
      write_address_data_log_force[4798] <= 6'h00;
      write_address_data_log_force[4799] <= 6'h00;
      write_address_data_log_force[4800] <= 6'h00;
      write_address_data_log_force[4801] <= 6'h00;
      write_address_data_log_force[4802] <= 6'h00;
      write_address_data_log_force[4803] <= 6'h00;
      write_address_data_log_force[4804] <= 6'h00;
      write_address_data_log_force[4805] <= 6'h00;
      write_address_data_log_force[4806] <= 6'h00;
      write_address_data_log_force[4807] <= 6'h00;
      write_address_data_log_force[4808] <= 6'h00;
      write_address_data_log_force[4809] <= 6'h00;
      write_address_data_log_force[4810] <= 6'h00;
      write_address_data_log_force[4811] <= 6'h00;
      write_address_data_log_force[4812] <= 6'h00;
      write_address_data_log_force[4813] <= 6'h00;
      write_address_data_log_force[4814] <= 6'h00;
      write_address_data_log_force[4815] <= 6'h00;
      write_address_data_log_force[4816] <= 6'h00;
      write_address_data_log_force[4817] <= 6'h00;
      write_address_data_log_force[4818] <= 6'h00;
      write_address_data_log_force[4819] <= 6'h00;
      write_address_data_log_force[4820] <= 6'h00;
      write_address_data_log_force[4821] <= 6'h00;
      write_address_data_log_force[4822] <= 6'h00;
      write_address_data_log_force[4823] <= 6'h00;
      write_address_data_log_force[4824] <= 6'h00;
      write_address_data_log_force[4825] <= 6'h00;
      write_address_data_log_force[4826] <= 6'h00;
      write_address_data_log_force[4827] <= 6'h00;
      write_address_data_log_force[4828] <= 6'h00;
      write_address_data_log_force[4829] <= 6'h00;
      write_address_data_log_force[4830] <= 6'h00;
      write_address_data_log_force[4831] <= 6'h00;
      write_address_data_log_force[4832] <= 6'h00;
      write_address_data_log_force[4833] <= 6'h00;
      write_address_data_log_force[4834] <= 6'h00;
      write_address_data_log_force[4835] <= 6'h00;
      write_address_data_log_force[4836] <= 6'h00;
      write_address_data_log_force[4837] <= 6'h00;
      write_address_data_log_force[4838] <= 6'h00;
      write_address_data_log_force[4839] <= 6'h00;
      write_address_data_log_force[4840] <= 6'h00;
      write_address_data_log_force[4841] <= 6'h00;
      write_address_data_log_force[4842] <= 6'h00;
      write_address_data_log_force[4843] <= 6'h00;
      write_address_data_log_force[4844] <= 6'h00;
      write_address_data_log_force[4845] <= 6'h00;
      write_address_data_log_force[4846] <= 6'h00;
      write_address_data_log_force[4847] <= 6'h00;
      write_address_data_log_force[4848] <= 6'h00;
      write_address_data_log_force[4849] <= 6'h00;
      write_address_data_log_force[4850] <= 6'h00;
      write_address_data_log_force[4851] <= 6'h00;
      write_address_data_log_force[4852] <= 6'h00;
      write_address_data_log_force[4853] <= 6'h00;
      write_address_data_log_force[4854] <= 6'h00;
      write_address_data_log_force[4855] <= 6'h00;
      write_address_data_log_force[4856] <= 6'h00;
      write_address_data_log_force[4857] <= 6'h00;
      write_address_data_log_force[4858] <= 6'h00;
      write_address_data_log_force[4859] <= 6'h00;
      write_address_data_log_force[4860] <= 6'h00;
      write_address_data_log_force[4861] <= 6'h00;
      write_address_data_log_force[4862] <= 6'h00;
      write_address_data_log_force[4863] <= 6'h00;
      write_address_data_log_force[4864] <= 6'h00;
      write_address_data_log_force[4865] <= 6'h00;
      write_address_data_log_force[4866] <= 6'h00;
      write_address_data_log_force[4867] <= 6'h00;
      write_address_data_log_force[4868] <= 6'h00;
      write_address_data_log_force[4869] <= 6'h00;
      write_address_data_log_force[4870] <= 6'h00;
      write_address_data_log_force[4871] <= 6'h00;
      write_address_data_log_force[4872] <= 6'h00;
      write_address_data_log_force[4873] <= 6'h00;
      write_address_data_log_force[4874] <= 6'h00;
      write_address_data_log_force[4875] <= 6'h00;
      write_address_data_log_force[4876] <= 6'h00;
      write_address_data_log_force[4877] <= 6'h00;
      write_address_data_log_force[4878] <= 6'h00;
      write_address_data_log_force[4879] <= 6'h00;
      write_address_data_log_force[4880] <= 6'h00;
      write_address_data_log_force[4881] <= 6'h00;
      write_address_data_log_force[4882] <= 6'h00;
      write_address_data_log_force[4883] <= 6'h00;
      write_address_data_log_force[4884] <= 6'h00;
      write_address_data_log_force[4885] <= 6'h00;
      write_address_data_log_force[4886] <= 6'h00;
      write_address_data_log_force[4887] <= 6'h00;
      write_address_data_log_force[4888] <= 6'h00;
      write_address_data_log_force[4889] <= 6'h00;
      write_address_data_log_force[4890] <= 6'h00;
      write_address_data_log_force[4891] <= 6'h00;
      write_address_data_log_force[4892] <= 6'h00;
      write_address_data_log_force[4893] <= 6'h00;
      write_address_data_log_force[4894] <= 6'h00;
      write_address_data_log_force[4895] <= 6'h00;
      write_address_data_log_force[4896] <= 6'h00;
      write_address_data_log_force[4897] <= 6'h00;
      write_address_data_log_force[4898] <= 6'h00;
      write_address_data_log_force[4899] <= 6'h00;
      write_address_data_log_force[4900] <= 6'h00;
      write_address_data_log_force[4901] <= 6'h00;
      write_address_data_log_force[4902] <= 6'h00;
      write_address_data_log_force[4903] <= 6'h00;
      write_address_data_log_force[4904] <= 6'h00;
      write_address_data_log_force[4905] <= 6'h00;
      write_address_data_log_force[4906] <= 6'h00;
      write_address_data_log_force[4907] <= 6'h00;
      write_address_data_log_force[4908] <= 6'h00;
      write_address_data_log_force[4909] <= 6'h00;
      write_address_data_log_force[4910] <= 6'h00;
      write_address_data_log_force[4911] <= 6'h00;
      write_address_data_log_force[4912] <= 6'h00;
      write_address_data_log_force[4913] <= 6'h00;
      write_address_data_log_force[4914] <= 6'h00;
      write_address_data_log_force[4915] <= 6'h00;
      write_address_data_log_force[4916] <= 6'h00;
      write_address_data_log_force[4917] <= 6'h00;
      write_address_data_log_force[4918] <= 6'h00;
      write_address_data_log_force[4919] <= 6'h00;
      write_address_data_log_force[4920] <= 6'h00;
      write_address_data_log_force[4921] <= 6'h00;
      write_address_data_log_force[4922] <= 6'h00;
      write_address_data_log_force[4923] <= 6'h00;
      write_address_data_log_force[4924] <= 6'h00;
      write_address_data_log_force[4925] <= 6'h00;
      write_address_data_log_force[4926] <= 6'h00;
      write_address_data_log_force[4927] <= 6'h00;
      write_address_data_log_force[4928] <= 6'h00;
      write_address_data_log_force[4929] <= 6'h00;
      write_address_data_log_force[4930] <= 6'h00;
      write_address_data_log_force[4931] <= 6'h00;
      write_address_data_log_force[4932] <= 6'h00;
      write_address_data_log_force[4933] <= 6'h00;
      write_address_data_log_force[4934] <= 6'h00;
      write_address_data_log_force[4935] <= 6'h00;
      write_address_data_log_force[4936] <= 6'h00;
      write_address_data_log_force[4937] <= 6'h00;
      write_address_data_log_force[4938] <= 6'h00;
      write_address_data_log_force[4939] <= 6'h00;
      write_address_data_log_force[4940] <= 6'h00;
      write_address_data_log_force[4941] <= 6'h00;
      write_address_data_log_force[4942] <= 6'h00;
      write_address_data_log_force[4943] <= 6'h00;
      write_address_data_log_force[4944] <= 6'h00;
      write_address_data_log_force[4945] <= 6'h00;
      write_address_data_log_force[4946] <= 6'h00;
      write_address_data_log_force[4947] <= 6'h00;
      write_address_data_log_force[4948] <= 6'h00;
      write_address_data_log_force[4949] <= 6'h00;
      write_address_data_log_force[4950] <= 6'h00;
      write_address_data_log_force[4951] <= 6'h00;
      write_address_data_log_force[4952] <= 6'h00;
      write_address_data_log_force[4953] <= 6'h00;
      write_address_data_log_force[4954] <= 6'h00;
      write_address_data_log_force[4955] <= 6'h00;
      write_address_data_log_force[4956] <= 6'h00;
      write_address_data_log_force[4957] <= 6'h00;
      write_address_data_log_force[4958] <= 6'h00;
      write_address_data_log_force[4959] <= 6'h00;
      write_address_data_log_force[4960] <= 6'h00;
      write_address_data_log_force[4961] <= 6'h00;
      write_address_data_log_force[4962] <= 6'h00;
      write_address_data_log_force[4963] <= 6'h00;
      write_address_data_log_force[4964] <= 6'h00;
      write_address_data_log_force[4965] <= 6'h00;
      write_address_data_log_force[4966] <= 6'h00;
      write_address_data_log_force[4967] <= 6'h00;
      write_address_data_log_force[4968] <= 6'h00;
      write_address_data_log_force[4969] <= 6'h00;
      write_address_data_log_force[4970] <= 6'h00;
      write_address_data_log_force[4971] <= 6'h00;
      write_address_data_log_force[4972] <= 6'h00;
      write_address_data_log_force[4973] <= 6'h00;
      write_address_data_log_force[4974] <= 6'h00;
      write_address_data_log_force[4975] <= 6'h00;
      write_address_data_log_force[4976] <= 6'h00;
      write_address_data_log_force[4977] <= 6'h00;
      write_address_data_log_force[4978] <= 6'h00;
      write_address_data_log_force[4979] <= 6'h00;
      write_address_data_log_force[4980] <= 6'h00;
      write_address_data_log_force[4981] <= 6'h00;
      write_address_data_log_force[4982] <= 6'h00;
      write_address_data_log_force[4983] <= 6'h00;
      write_address_data_log_force[4984] <= 6'h00;
      write_address_data_log_force[4985] <= 6'h00;
      write_address_data_log_force[4986] <= 6'h00;
      write_address_data_log_force[4987] <= 6'h00;
      write_address_data_log_force[4988] <= 6'h00;
      write_address_data_log_force[4989] <= 6'h00;
      write_address_data_log_force[4990] <= 6'h00;
      write_address_data_log_force[4991] <= 6'h00;
      write_address_data_log_force[4992] <= 6'h00;
      write_address_data_log_force[4993] <= 6'h00;
      write_address_data_log_force[4994] <= 6'h00;
      write_address_data_log_force[4995] <= 6'h00;
      write_address_data_log_force[4996] <= 6'h00;
      write_address_data_log_force[4997] <= 6'h00;
      write_address_data_log_force[4998] <= 6'h00;
      write_address_data_log_force[4999] <= 6'h00;
      write_address_data_log_force[5000] <= 6'h00;
      write_address_data_log_force[5001] <= 6'h00;
      write_address_data_log_force[5002] <= 6'h00;
      write_address_data_log_force[5003] <= 6'h00;
      write_address_data_log_force[5004] <= 6'h00;
      write_address_data_log_force[5005] <= 6'h00;
      write_address_data_log_force[5006] <= 6'h00;
      write_address_data_log_force[5007] <= 6'h00;
      write_address_data_log_force[5008] <= 6'h00;
      write_address_data_log_force[5009] <= 6'h00;
      write_address_data_log_force[5010] <= 6'h00;
      write_address_data_log_force[5011] <= 6'h00;
      write_address_data_log_force[5012] <= 6'h00;
      write_address_data_log_force[5013] <= 6'h00;
      write_address_data_log_force[5014] <= 6'h00;
      write_address_data_log_force[5015] <= 6'h00;
      write_address_data_log_force[5016] <= 6'h00;
      write_address_data_log_force[5017] <= 6'h00;
      write_address_data_log_force[5018] <= 6'h00;
      write_address_data_log_force[5019] <= 6'h00;
      write_address_data_log_force[5020] <= 6'h00;
      write_address_data_log_force[5021] <= 6'h00;
      write_address_data_log_force[5022] <= 6'h00;
      write_address_data_log_force[5023] <= 6'h00;
      write_address_data_log_force[5024] <= 6'h00;
      write_address_data_log_force[5025] <= 6'h00;
      write_address_data_log_force[5026] <= 6'h00;
      write_address_data_log_force[5027] <= 6'h00;
      write_address_data_log_force[5028] <= 6'h00;
      write_address_data_log_force[5029] <= 6'h00;
      write_address_data_log_force[5030] <= 6'h00;
      write_address_data_log_force[5031] <= 6'h00;
      write_address_data_log_force[5032] <= 6'h00;
      write_address_data_log_force[5033] <= 6'h00;
      write_address_data_log_force[5034] <= 6'h00;
      write_address_data_log_force[5035] <= 6'h00;
      write_address_data_log_force[5036] <= 6'h00;
      write_address_data_log_force[5037] <= 6'h00;
      write_address_data_log_force[5038] <= 6'h00;
      write_address_data_log_force[5039] <= 6'h00;
      write_address_data_log_force[5040] <= 6'h00;
      write_address_data_log_force[5041] <= 6'h00;
      write_address_data_log_force[5042] <= 6'h00;
      write_address_data_log_force[5043] <= 6'h00;
      write_address_data_log_force[5044] <= 6'h00;
      write_address_data_log_force[5045] <= 6'h00;
      write_address_data_log_force[5046] <= 6'h00;
      write_address_data_log_force[5047] <= 6'h00;
      write_address_data_log_force[5048] <= 6'h00;
      write_address_data_log_force[5049] <= 6'h00;
      write_address_data_log_force[5050] <= 6'h00;
      write_address_data_log_force[5051] <= 6'h00;
      write_address_data_log_force[5052] <= 6'h00;
      write_address_data_log_force[5053] <= 6'h00;
      write_address_data_log_force[5054] <= 6'h00;
      write_address_data_log_force[5055] <= 6'h00;
      write_address_data_log_force[5056] <= 6'h00;
      write_address_data_log_force[5057] <= 6'h00;
      write_address_data_log_force[5058] <= 6'h00;
      write_address_data_log_force[5059] <= 6'h00;
      write_address_data_log_force[5060] <= 6'h00;
      write_address_data_log_force[5061] <= 6'h00;
      write_address_data_log_force[5062] <= 6'h00;
      write_address_data_log_force[5063] <= 6'h00;
      write_address_data_log_force[5064] <= 6'h00;
      write_address_data_log_force[5065] <= 6'h00;
      write_address_data_log_force[5066] <= 6'h00;
      write_address_data_log_force[5067] <= 6'h00;
      write_address_data_log_force[5068] <= 6'h00;
      write_address_data_log_force[5069] <= 6'h00;
      write_address_data_log_force[5070] <= 6'h00;
      write_address_data_log_force[5071] <= 6'h00;
      write_address_data_log_force[5072] <= 6'h00;
      write_address_data_log_force[5073] <= 6'h00;
      write_address_data_log_force[5074] <= 6'h00;
      write_address_data_log_force[5075] <= 6'h00;
      write_address_data_log_force[5076] <= 6'h00;
      write_address_data_log_force[5077] <= 6'h00;
      write_address_data_log_force[5078] <= 6'h00;
      write_address_data_log_force[5079] <= 6'h00;
      write_address_data_log_force[5080] <= 6'h00;
      write_address_data_log_force[5081] <= 6'h00;
      write_address_data_log_force[5082] <= 6'h00;
      write_address_data_log_force[5083] <= 6'h00;
      write_address_data_log_force[5084] <= 6'h00;
      write_address_data_log_force[5085] <= 6'h00;
      write_address_data_log_force[5086] <= 6'h00;
      write_address_data_log_force[5087] <= 6'h00;
      write_address_data_log_force[5088] <= 6'h00;
      write_address_data_log_force[5089] <= 6'h00;
      write_address_data_log_force[5090] <= 6'h00;
      write_address_data_log_force[5091] <= 6'h00;
      write_address_data_log_force[5092] <= 6'h00;
      write_address_data_log_force[5093] <= 6'h00;
      write_address_data_log_force[5094] <= 6'h00;
      write_address_data_log_force[5095] <= 6'h00;
      write_address_data_log_force[5096] <= 6'h00;
      write_address_data_log_force[5097] <= 6'h00;
      write_address_data_log_force[5098] <= 6'h00;
      write_address_data_log_force[5099] <= 6'h00;
      write_address_data_log_force[5100] <= 6'h00;
      write_address_data_log_force[5101] <= 6'h00;
      write_address_data_log_force[5102] <= 6'h00;
      write_address_data_log_force[5103] <= 6'h00;
      write_address_data_log_force[5104] <= 6'h00;
      write_address_data_log_force[5105] <= 6'h00;
      write_address_data_log_force[5106] <= 6'h00;
      write_address_data_log_force[5107] <= 6'h00;
      write_address_data_log_force[5108] <= 6'h00;
      write_address_data_log_force[5109] <= 6'h00;
      write_address_data_log_force[5110] <= 6'h00;
      write_address_data_log_force[5111] <= 6'h00;
      write_address_data_log_force[5112] <= 6'h00;
      write_address_data_log_force[5113] <= 6'h00;
      write_address_data_log_force[5114] <= 6'h00;
      write_address_data_log_force[5115] <= 6'h00;
      write_address_data_log_force[5116] <= 6'h00;
      write_address_data_log_force[5117] <= 6'h00;
      write_address_data_log_force[5118] <= 6'h00;
      write_address_data_log_force[5119] <= 6'h00;
      write_address_data_log_force[5120] <= 6'h00;
      write_address_data_log_force[5121] <= 6'h00;
      write_address_data_log_force[5122] <= 6'h00;
      write_address_data_log_force[5123] <= 6'h00;
      write_address_data_log_force[5124] <= 6'h00;
      write_address_data_log_force[5125] <= 6'h00;
      write_address_data_log_force[5126] <= 6'h00;
      write_address_data_log_force[5127] <= 6'h00;
      write_address_data_log_force[5128] <= 6'h00;
      write_address_data_log_force[5129] <= 6'h00;
      write_address_data_log_force[5130] <= 6'h00;
      write_address_data_log_force[5131] <= 6'h00;
      write_address_data_log_force[5132] <= 6'h00;
      write_address_data_log_force[5133] <= 6'h00;
      write_address_data_log_force[5134] <= 6'h00;
      write_address_data_log_force[5135] <= 6'h00;
      write_address_data_log_force[5136] <= 6'h00;
      write_address_data_log_force[5137] <= 6'h00;
      write_address_data_log_force[5138] <= 6'h00;
      write_address_data_log_force[5139] <= 6'h00;
      write_address_data_log_force[5140] <= 6'h00;
      write_address_data_log_force[5141] <= 6'h00;
      write_address_data_log_force[5142] <= 6'h00;
      write_address_data_log_force[5143] <= 6'h00;
      write_address_data_log_force[5144] <= 6'h00;
      write_address_data_log_force[5145] <= 6'h00;
      write_address_data_log_force[5146] <= 6'h00;
      write_address_data_log_force[5147] <= 6'h00;
      write_address_data_log_force[5148] <= 6'h00;
      write_address_data_log_force[5149] <= 6'h00;
      write_address_data_log_force[5150] <= 6'h00;
      write_address_data_log_force[5151] <= 6'h00;
      write_address_data_log_force[5152] <= 6'h00;
      write_address_data_log_force[5153] <= 6'h00;
      write_address_data_log_force[5154] <= 6'h00;
      write_address_data_log_force[5155] <= 6'h00;
      write_address_data_log_force[5156] <= 6'h00;
      write_address_data_log_force[5157] <= 6'h00;
      write_address_data_log_force[5158] <= 6'h00;
      write_address_data_log_force[5159] <= 6'h00;
      write_address_data_log_force[5160] <= 6'h00;
      write_address_data_log_force[5161] <= 6'h00;
      write_address_data_log_force[5162] <= 6'h00;
      write_address_data_log_force[5163] <= 6'h00;
      write_address_data_log_force[5164] <= 6'h00;
      write_address_data_log_force[5165] <= 6'h00;
      write_address_data_log_force[5166] <= 6'h00;
      write_address_data_log_force[5167] <= 6'h00;
      write_address_data_log_force[5168] <= 6'h00;
      write_address_data_log_force[5169] <= 6'h00;
      write_address_data_log_force[5170] <= 6'h00;
      write_address_data_log_force[5171] <= 6'h00;
      write_address_data_log_force[5172] <= 6'h00;
      write_address_data_log_force[5173] <= 6'h00;
      write_address_data_log_force[5174] <= 6'h00;
      write_address_data_log_force[5175] <= 6'h00;
      write_address_data_log_force[5176] <= 6'h00;
      write_address_data_log_force[5177] <= 6'h00;
      write_address_data_log_force[5178] <= 6'h00;
      write_address_data_log_force[5179] <= 6'h00;
      write_address_data_log_force[5180] <= 6'h00;
      write_address_data_log_force[5181] <= 6'h00;
      write_address_data_log_force[5182] <= 6'h00;
      write_address_data_log_force[5183] <= 6'h00;
      write_address_data_log_force[5184] <= 6'h00;
      write_address_data_log_force[5185] <= 6'h00;
      write_address_data_log_force[5186] <= 6'h00;
      write_address_data_log_force[5187] <= 6'h00;
      write_address_data_log_force[5188] <= 6'h00;
      write_address_data_log_force[5189] <= 6'h00;
      write_address_data_log_force[5190] <= 6'h00;
      write_address_data_log_force[5191] <= 6'h00;
      write_address_data_log_force[5192] <= 6'h00;
      write_address_data_log_force[5193] <= 6'h00;
      write_address_data_log_force[5194] <= 6'h00;
      write_address_data_log_force[5195] <= 6'h00;
      write_address_data_log_force[5196] <= 6'h00;
      write_address_data_log_force[5197] <= 6'h00;
      write_address_data_log_force[5198] <= 6'h00;
      write_address_data_log_force[5199] <= 6'h00;
      write_address_data_log_force[5200] <= 6'h00;
      write_address_data_log_force[5201] <= 6'h00;
      write_address_data_log_force[5202] <= 6'h00;
      write_address_data_log_force[5203] <= 6'h00;
      write_address_data_log_force[5204] <= 6'h00;
      write_address_data_log_force[5205] <= 6'h00;
      write_address_data_log_force[5206] <= 6'h00;
      write_address_data_log_force[5207] <= 6'h00;
      write_address_data_log_force[5208] <= 6'h00;
      write_address_data_log_force[5209] <= 6'h00;
      write_address_data_log_force[5210] <= 6'h00;
      write_address_data_log_force[5211] <= 6'h00;
      write_address_data_log_force[5212] <= 6'h00;
      write_address_data_log_force[5213] <= 6'h00;
      write_address_data_log_force[5214] <= 6'h00;
      write_address_data_log_force[5215] <= 6'h00;
      write_address_data_log_force[5216] <= 6'h00;
      write_address_data_log_force[5217] <= 6'h00;
      write_address_data_log_force[5218] <= 6'h00;
      write_address_data_log_force[5219] <= 6'h00;
      write_address_data_log_force[5220] <= 6'h00;
      write_address_data_log_force[5221] <= 6'h00;
      write_address_data_log_force[5222] <= 6'h00;
      write_address_data_log_force[5223] <= 6'h00;
      write_address_data_log_force[5224] <= 6'h00;
      write_address_data_log_force[5225] <= 6'h00;
      write_address_data_log_force[5226] <= 6'h00;
      write_address_data_log_force[5227] <= 6'h00;
      write_address_data_log_force[5228] <= 6'h00;
      write_address_data_log_force[5229] <= 6'h00;
      write_address_data_log_force[5230] <= 6'h00;
      write_address_data_log_force[5231] <= 6'h00;
      write_address_data_log_force[5232] <= 6'h00;
      write_address_data_log_force[5233] <= 6'h00;
      write_address_data_log_force[5234] <= 6'h00;
      write_address_data_log_force[5235] <= 6'h00;
      write_address_data_log_force[5236] <= 6'h00;
      write_address_data_log_force[5237] <= 6'h00;
      write_address_data_log_force[5238] <= 6'h00;
      write_address_data_log_force[5239] <= 6'h00;
      write_address_data_log_force[5240] <= 6'h00;
      write_address_data_log_force[5241] <= 6'h00;
      write_address_data_log_force[5242] <= 6'h00;
      write_address_data_log_force[5243] <= 6'h00;
      write_address_data_log_force[5244] <= 6'h00;
      write_address_data_log_force[5245] <= 6'h00;
      write_address_data_log_force[5246] <= 6'h00;
      write_address_data_log_force[5247] <= 6'h00;
      write_address_data_log_force[5248] <= 6'h00;
      write_address_data_log_force[5249] <= 6'h00;
      write_address_data_log_force[5250] <= 6'h00;
      write_address_data_log_force[5251] <= 6'h00;
      write_address_data_log_force[5252] <= 6'h00;
      write_address_data_log_force[5253] <= 6'h00;
      write_address_data_log_force[5254] <= 6'h00;
      write_address_data_log_force[5255] <= 6'h00;
      write_address_data_log_force[5256] <= 6'h00;
      write_address_data_log_force[5257] <= 6'h00;
      write_address_data_log_force[5258] <= 6'h00;
      write_address_data_log_force[5259] <= 6'h00;
      write_address_data_log_force[5260] <= 6'h00;
      write_address_data_log_force[5261] <= 6'h00;
      write_address_data_log_force[5262] <= 6'h00;
      write_address_data_log_force[5263] <= 6'h00;
      write_address_data_log_force[5264] <= 6'h00;
      write_address_data_log_force[5265] <= 6'h00;
      write_address_data_log_force[5266] <= 6'h00;
      write_address_data_log_force[5267] <= 6'h00;
      write_address_data_log_force[5268] <= 6'h00;
      write_address_data_log_force[5269] <= 6'h00;
      write_address_data_log_force[5270] <= 6'h00;
      write_address_data_log_force[5271] <= 6'h00;
      write_address_data_log_force[5272] <= 6'h00;
      write_address_data_log_force[5273] <= 6'h00;
      write_address_data_log_force[5274] <= 6'h00;
      write_address_data_log_force[5275] <= 6'h00;
      write_address_data_log_force[5276] <= 6'h00;
      write_address_data_log_force[5277] <= 6'h00;
      write_address_data_log_force[5278] <= 6'h00;
      write_address_data_log_force[5279] <= 6'h00;
      write_address_data_log_force[5280] <= 6'h00;
      write_address_data_log_force[5281] <= 6'h00;
      write_address_data_log_force[5282] <= 6'h00;
      write_address_data_log_force[5283] <= 6'h00;
      write_address_data_log_force[5284] <= 6'h00;
      write_address_data_log_force[5285] <= 6'h00;
      write_address_data_log_force[5286] <= 6'h00;
      write_address_data_log_force[5287] <= 6'h00;
      write_address_data_log_force[5288] <= 6'h00;
      write_address_data_log_force[5289] <= 6'h00;
      write_address_data_log_force[5290] <= 6'h00;
      write_address_data_log_force[5291] <= 6'h00;
      write_address_data_log_force[5292] <= 6'h00;
      write_address_data_log_force[5293] <= 6'h00;
      write_address_data_log_force[5294] <= 6'h00;
      write_address_data_log_force[5295] <= 6'h00;
      write_address_data_log_force[5296] <= 6'h00;
      write_address_data_log_force[5297] <= 6'h00;
      write_address_data_log_force[5298] <= 6'h00;
      write_address_data_log_force[5299] <= 6'h00;
      write_address_data_log_force[5300] <= 6'h00;
      write_address_data_log_force[5301] <= 6'h00;
      write_address_data_log_force[5302] <= 6'h00;
      write_address_data_log_force[5303] <= 6'h00;
      write_address_data_log_force[5304] <= 6'h00;
      write_address_data_log_force[5305] <= 6'h00;
      write_address_data_log_force[5306] <= 6'h00;
      write_address_data_log_force[5307] <= 6'h00;
      write_address_data_log_force[5308] <= 6'h00;
      write_address_data_log_force[5309] <= 6'h00;
      write_address_data_log_force[5310] <= 6'h00;
      write_address_data_log_force[5311] <= 6'h00;
      write_address_data_log_force[5312] <= 6'h00;
      write_address_data_log_force[5313] <= 6'h00;
      write_address_data_log_force[5314] <= 6'h00;
      write_address_data_log_force[5315] <= 6'h00;
      write_address_data_log_force[5316] <= 6'h00;
      write_address_data_log_force[5317] <= 6'h00;
      write_address_data_log_force[5318] <= 6'h00;
      write_address_data_log_force[5319] <= 6'h00;
      write_address_data_log_force[5320] <= 6'h00;
      write_address_data_log_force[5321] <= 6'h00;
      write_address_data_log_force[5322] <= 6'h00;
      write_address_data_log_force[5323] <= 6'h00;
      write_address_data_log_force[5324] <= 6'h00;
      write_address_data_log_force[5325] <= 6'h00;
      write_address_data_log_force[5326] <= 6'h00;
      write_address_data_log_force[5327] <= 6'h00;
      write_address_data_log_force[5328] <= 6'h00;
      write_address_data_log_force[5329] <= 6'h00;
      write_address_data_log_force[5330] <= 6'h00;
      write_address_data_log_force[5331] <= 6'h00;
      write_address_data_log_force[5332] <= 6'h00;
      write_address_data_log_force[5333] <= 6'h00;
      write_address_data_log_force[5334] <= 6'h00;
      write_address_data_log_force[5335] <= 6'h00;
      write_address_data_log_force[5336] <= 6'h00;
      write_address_data_log_force[5337] <= 6'h00;
      write_address_data_log_force[5338] <= 6'h00;
      write_address_data_log_force[5339] <= 6'h00;
      write_address_data_log_force[5340] <= 6'h00;
      write_address_data_log_force[5341] <= 6'h00;
      write_address_data_log_force[5342] <= 6'h00;
      write_address_data_log_force[5343] <= 6'h00;
      write_address_data_log_force[5344] <= 6'h00;
      write_address_data_log_force[5345] <= 6'h00;
      write_address_data_log_force[5346] <= 6'h00;
      write_address_data_log_force[5347] <= 6'h00;
      write_address_data_log_force[5348] <= 6'h00;
      write_address_data_log_force[5349] <= 6'h00;
      write_address_data_log_force[5350] <= 6'h00;
      write_address_data_log_force[5351] <= 6'h00;
      write_address_data_log_force[5352] <= 6'h00;
      write_address_data_log_force[5353] <= 6'h00;
      write_address_data_log_force[5354] <= 6'h00;
      write_address_data_log_force[5355] <= 6'h00;
      write_address_data_log_force[5356] <= 6'h00;
      write_address_data_log_force[5357] <= 6'h00;
      write_address_data_log_force[5358] <= 6'h00;
      write_address_data_log_force[5359] <= 6'h00;
      write_address_data_log_force[5360] <= 6'h00;
      write_address_data_log_force[5361] <= 6'h00;
      write_address_data_log_force[5362] <= 6'h00;
      write_address_data_log_force[5363] <= 6'h00;
      write_address_data_log_force[5364] <= 6'h00;
      write_address_data_log_force[5365] <= 6'h00;
      write_address_data_log_force[5366] <= 6'h00;
      write_address_data_log_force[5367] <= 6'h00;
      write_address_data_log_force[5368] <= 6'h00;
      write_address_data_log_force[5369] <= 6'h00;
      write_address_data_log_force[5370] <= 6'h00;
      write_address_data_log_force[5371] <= 6'h00;
      write_address_data_log_force[5372] <= 6'h00;
      write_address_data_log_force[5373] <= 6'h00;
      write_address_data_log_force[5374] <= 6'h00;
      write_address_data_log_force[5375] <= 6'h00;
      write_address_data_log_force[5376] <= 6'h00;
      write_address_data_log_force[5377] <= 6'h00;
      write_address_data_log_force[5378] <= 6'h00;
      write_address_data_log_force[5379] <= 6'h00;
      write_address_data_log_force[5380] <= 6'h00;
      write_address_data_log_force[5381] <= 6'h00;
      write_address_data_log_force[5382] <= 6'h00;
      write_address_data_log_force[5383] <= 6'h00;
      write_address_data_log_force[5384] <= 6'h00;
      write_address_data_log_force[5385] <= 6'h00;
      write_address_data_log_force[5386] <= 6'h00;
      write_address_data_log_force[5387] <= 6'h00;
      write_address_data_log_force[5388] <= 6'h00;
      write_address_data_log_force[5389] <= 6'h00;
      write_address_data_log_force[5390] <= 6'h00;
      write_address_data_log_force[5391] <= 6'h00;
      write_address_data_log_force[5392] <= 6'h00;
      write_address_data_log_force[5393] <= 6'h00;
      write_address_data_log_force[5394] <= 6'h00;
      write_address_data_log_force[5395] <= 6'h00;
      write_address_data_log_force[5396] <= 6'h00;
      write_address_data_log_force[5397] <= 6'h00;
      write_address_data_log_force[5398] <= 6'h00;
      write_address_data_log_force[5399] <= 6'h00;
      write_address_data_log_force[5400] <= 6'h00;
      write_address_data_log_force[5401] <= 6'h00;
      write_address_data_log_force[5402] <= 6'h00;
      write_address_data_log_force[5403] <= 6'h00;
      write_address_data_log_force[5404] <= 6'h00;
      write_address_data_log_force[5405] <= 6'h00;
      write_address_data_log_force[5406] <= 6'h00;
      write_address_data_log_force[5407] <= 6'h00;
      write_address_data_log_force[5408] <= 6'h00;
      write_address_data_log_force[5409] <= 6'h00;
      write_address_data_log_force[5410] <= 6'h00;
      write_address_data_log_force[5411] <= 6'h00;
      write_address_data_log_force[5412] <= 6'h00;
      write_address_data_log_force[5413] <= 6'h00;
      write_address_data_log_force[5414] <= 6'h00;
      write_address_data_log_force[5415] <= 6'h00;
      write_address_data_log_force[5416] <= 6'h00;
      write_address_data_log_force[5417] <= 6'h00;
      write_address_data_log_force[5418] <= 6'h00;
      write_address_data_log_force[5419] <= 6'h00;
      write_address_data_log_force[5420] <= 6'h00;
      write_address_data_log_force[5421] <= 6'h00;
      write_address_data_log_force[5422] <= 6'h00;
      write_address_data_log_force[5423] <= 6'h00;
      write_address_data_log_force[5424] <= 6'h00;
      write_address_data_log_force[5425] <= 6'h00;
      write_address_data_log_force[5426] <= 6'h00;
      write_address_data_log_force[5427] <= 6'h00;
      write_address_data_log_force[5428] <= 6'h00;
      write_address_data_log_force[5429] <= 6'h00;
      write_address_data_log_force[5430] <= 6'h00;
      write_address_data_log_force[5431] <= 6'h00;
      write_address_data_log_force[5432] <= 6'h00;
      write_address_data_log_force[5433] <= 6'h00;
      write_address_data_log_force[5434] <= 6'h00;
      write_address_data_log_force[5435] <= 6'h00;
      write_address_data_log_force[5436] <= 6'h00;
      write_address_data_log_force[5437] <= 6'h00;
      write_address_data_log_force[5438] <= 6'h00;
      write_address_data_log_force[5439] <= 6'h00;
      write_address_data_log_force[5440] <= 6'h00;
      write_address_data_log_force[5441] <= 6'h00;
      write_address_data_log_force[5442] <= 6'h00;
      write_address_data_log_force[5443] <= 6'h00;
      write_address_data_log_force[5444] <= 6'h00;
      write_address_data_log_force[5445] <= 6'h00;
      write_address_data_log_force[5446] <= 6'h00;
      write_address_data_log_force[5447] <= 6'h00;
      write_address_data_log_force[5448] <= 6'h00;
      write_address_data_log_force[5449] <= 6'h00;
      write_address_data_log_force[5450] <= 6'h00;
      write_address_data_log_force[5451] <= 6'h00;
      write_address_data_log_force[5452] <= 6'h00;
      write_address_data_log_force[5453] <= 6'h00;
      write_address_data_log_force[5454] <= 6'h00;
      write_address_data_log_force[5455] <= 6'h00;
      write_address_data_log_force[5456] <= 6'h00;
      write_address_data_log_force[5457] <= 6'h00;
      write_address_data_log_force[5458] <= 6'h00;
      write_address_data_log_force[5459] <= 6'h00;
      write_address_data_log_force[5460] <= 6'h00;
      write_address_data_log_force[5461] <= 6'h00;
      write_address_data_log_force[5462] <= 6'h00;
      write_address_data_log_force[5463] <= 6'h00;
      write_address_data_log_force[5464] <= 6'h00;
      write_address_data_log_force[5465] <= 6'h00;
      write_address_data_log_force[5466] <= 6'h00;
      write_address_data_log_force[5467] <= 6'h00;
      write_address_data_log_force[5468] <= 6'h00;
      write_address_data_log_force[5469] <= 6'h00;
      write_address_data_log_force[5470] <= 6'h00;
      write_address_data_log_force[5471] <= 6'h00;
      write_address_data_log_force[5472] <= 6'h00;
      write_address_data_log_force[5473] <= 6'h00;
      write_address_data_log_force[5474] <= 6'h00;
      write_address_data_log_force[5475] <= 6'h00;
      write_address_data_log_force[5476] <= 6'h00;
      write_address_data_log_force[5477] <= 6'h00;
      write_address_data_log_force[5478] <= 6'h00;
      write_address_data_log_force[5479] <= 6'h00;
      write_address_data_log_force[5480] <= 6'h00;
      write_address_data_log_force[5481] <= 6'h00;
      write_address_data_log_force[5482] <= 6'h00;
      write_address_data_log_force[5483] <= 6'h00;
      write_address_data_log_force[5484] <= 6'h00;
      write_address_data_log_force[5485] <= 6'h00;
      write_address_data_log_force[5486] <= 6'h00;
      write_address_data_log_force[5487] <= 6'h00;
      write_address_data_log_force[5488] <= 6'h00;
      write_address_data_log_force[5489] <= 6'h00;
      write_address_data_log_force[5490] <= 6'h00;
      write_address_data_log_force[5491] <= 6'h00;
      write_address_data_log_force[5492] <= 6'h00;
      write_address_data_log_force[5493] <= 6'h00;
      write_address_data_log_force[5494] <= 6'h00;
      write_address_data_log_force[5495] <= 6'h00;
      write_address_data_log_force[5496] <= 6'h00;
      write_address_data_log_force[5497] <= 6'h00;
      write_address_data_log_force[5498] <= 6'h00;
      write_address_data_log_force[5499] <= 6'h00;
      write_address_data_log_force[5500] <= 6'h00;
      write_address_data_log_force[5501] <= 6'h00;
      write_address_data_log_force[5502] <= 6'h00;
      write_address_data_log_force[5503] <= 6'h00;
      write_address_data_log_force[5504] <= 6'h00;
      write_address_data_log_force[5505] <= 6'h00;
      write_address_data_log_force[5506] <= 6'h00;
      write_address_data_log_force[5507] <= 6'h00;
      write_address_data_log_force[5508] <= 6'h00;
      write_address_data_log_force[5509] <= 6'h00;
      write_address_data_log_force[5510] <= 6'h00;
      write_address_data_log_force[5511] <= 6'h00;
      write_address_data_log_force[5512] <= 6'h00;
      write_address_data_log_force[5513] <= 6'h00;
      write_address_data_log_force[5514] <= 6'h00;
      write_address_data_log_force[5515] <= 6'h00;
      write_address_data_log_force[5516] <= 6'h00;
      write_address_data_log_force[5517] <= 6'h00;
      write_address_data_log_force[5518] <= 6'h00;
      write_address_data_log_force[5519] <= 6'h00;
      write_address_data_log_force[5520] <= 6'h00;
      write_address_data_log_force[5521] <= 6'h00;
      write_address_data_log_force[5522] <= 6'h00;
      write_address_data_log_force[5523] <= 6'h00;
      write_address_data_log_force[5524] <= 6'h00;
      write_address_data_log_force[5525] <= 6'h00;
      write_address_data_log_force[5526] <= 6'h00;
      write_address_data_log_force[5527] <= 6'h00;
      write_address_data_log_force[5528] <= 6'h00;
      write_address_data_log_force[5529] <= 6'h00;
      write_address_data_log_force[5530] <= 6'h00;
      write_address_data_log_force[5531] <= 6'h00;
      write_address_data_log_force[5532] <= 6'h00;
      write_address_data_log_force[5533] <= 6'h00;
      write_address_data_log_force[5534] <= 6'h00;
      write_address_data_log_force[5535] <= 6'h00;
      write_address_data_log_force[5536] <= 6'h00;
      write_address_data_log_force[5537] <= 6'h00;
      write_address_data_log_force[5538] <= 6'h00;
      write_address_data_log_force[5539] <= 6'h00;
      write_address_data_log_force[5540] <= 6'h00;
      write_address_data_log_force[5541] <= 6'h00;
      write_address_data_log_force[5542] <= 6'h00;
      write_address_data_log_force[5543] <= 6'h00;
      write_address_data_log_force[5544] <= 6'h00;
      write_address_data_log_force[5545] <= 6'h00;
      write_address_data_log_force[5546] <= 6'h00;
      write_address_data_log_force[5547] <= 6'h00;
      write_address_data_log_force[5548] <= 6'h00;
      write_address_data_log_force[5549] <= 6'h00;
      write_address_data_log_force[5550] <= 6'h00;
      write_address_data_log_force[5551] <= 6'h00;
      write_address_data_log_force[5552] <= 6'h00;
      write_address_data_log_force[5553] <= 6'h00;
      write_address_data_log_force[5554] <= 6'h00;
      write_address_data_log_force[5555] <= 6'h00;
      write_address_data_log_force[5556] <= 6'h00;
      write_address_data_log_force[5557] <= 6'h00;
      write_address_data_log_force[5558] <= 6'h00;
      write_address_data_log_force[5559] <= 6'h00;
      write_address_data_log_force[5560] <= 6'h00;
      write_address_data_log_force[5561] <= 6'h00;
      write_address_data_log_force[5562] <= 6'h00;
      write_address_data_log_force[5563] <= 6'h00;
      write_address_data_log_force[5564] <= 6'h00;
      write_address_data_log_force[5565] <= 6'h00;
      write_address_data_log_force[5566] <= 6'h00;
      write_address_data_log_force[5567] <= 6'h00;
      write_address_data_log_force[5568] <= 6'h00;
      write_address_data_log_force[5569] <= 6'h00;
      write_address_data_log_force[5570] <= 6'h00;
      write_address_data_log_force[5571] <= 6'h00;
      write_address_data_log_force[5572] <= 6'h00;
      write_address_data_log_force[5573] <= 6'h00;
      write_address_data_log_force[5574] <= 6'h00;
      write_address_data_log_force[5575] <= 6'h00;
      write_address_data_log_force[5576] <= 6'h00;
      write_address_data_log_force[5577] <= 6'h00;
      write_address_data_log_force[5578] <= 6'h00;
      write_address_data_log_force[5579] <= 6'h00;
      write_address_data_log_force[5580] <= 6'h00;
      write_address_data_log_force[5581] <= 6'h00;
      write_address_data_log_force[5582] <= 6'h00;
      write_address_data_log_force[5583] <= 6'h00;
      write_address_data_log_force[5584] <= 6'h00;
      write_address_data_log_force[5585] <= 6'h00;
      write_address_data_log_force[5586] <= 6'h00;
      write_address_data_log_force[5587] <= 6'h00;
      write_address_data_log_force[5588] <= 6'h00;
      write_address_data_log_force[5589] <= 6'h00;
      write_address_data_log_force[5590] <= 6'h00;
      write_address_data_log_force[5591] <= 6'h00;
      write_address_data_log_force[5592] <= 6'h00;
      write_address_data_log_force[5593] <= 6'h00;
      write_address_data_log_force[5594] <= 6'h00;
      write_address_data_log_force[5595] <= 6'h00;
      write_address_data_log_force[5596] <= 6'h00;
      write_address_data_log_force[5597] <= 6'h00;
      write_address_data_log_force[5598] <= 6'h00;
      write_address_data_log_force[5599] <= 6'h00;
      write_address_data_log_force[5600] <= 6'h00;
      write_address_data_log_force[5601] <= 6'h00;
      write_address_data_log_force[5602] <= 6'h00;
      write_address_data_log_force[5603] <= 6'h00;
      write_address_data_log_force[5604] <= 6'h00;
      write_address_data_log_force[5605] <= 6'h00;
      write_address_data_log_force[5606] <= 6'h00;
      write_address_data_log_force[5607] <= 6'h00;
      write_address_data_log_force[5608] <= 6'h00;
      write_address_data_log_force[5609] <= 6'h00;
      write_address_data_log_force[5610] <= 6'h00;
      write_address_data_log_force[5611] <= 6'h00;
      write_address_data_log_force[5612] <= 6'h00;
      write_address_data_log_force[5613] <= 6'h00;
      write_address_data_log_force[5614] <= 6'h00;
      write_address_data_log_force[5615] <= 6'h00;
      write_address_data_log_force[5616] <= 6'h00;
      write_address_data_log_force[5617] <= 6'h00;
      write_address_data_log_force[5618] <= 6'h00;
      write_address_data_log_force[5619] <= 6'h00;
      write_address_data_log_force[5620] <= 6'h00;
      write_address_data_log_force[5621] <= 6'h00;
      write_address_data_log_force[5622] <= 6'h00;
      write_address_data_log_force[5623] <= 6'h00;
      write_address_data_log_force[5624] <= 6'h00;
      write_address_data_log_force[5625] <= 6'h00;
      write_address_data_log_force[5626] <= 6'h00;
      write_address_data_log_force[5627] <= 6'h00;
      write_address_data_log_force[5628] <= 6'h00;
      write_address_data_log_force[5629] <= 6'h00;
      write_address_data_log_force[5630] <= 6'h00;
      write_address_data_log_force[5631] <= 6'h00;
      write_address_data_log_force[5632] <= 6'h00;
      write_address_data_log_force[5633] <= 6'h00;
      write_address_data_log_force[5634] <= 6'h00;
      write_address_data_log_force[5635] <= 6'h00;
      write_address_data_log_force[5636] <= 6'h00;
      write_address_data_log_force[5637] <= 6'h00;
      write_address_data_log_force[5638] <= 6'h00;
      write_address_data_log_force[5639] <= 6'h00;
      write_address_data_log_force[5640] <= 6'h00;
      write_address_data_log_force[5641] <= 6'h00;
      write_address_data_log_force[5642] <= 6'h00;
      write_address_data_log_force[5643] <= 6'h00;
      write_address_data_log_force[5644] <= 6'h00;
      write_address_data_log_force[5645] <= 6'h00;
      write_address_data_log_force[5646] <= 6'h00;
      write_address_data_log_force[5647] <= 6'h00;
      write_address_data_log_force[5648] <= 6'h00;
      write_address_data_log_force[5649] <= 6'h00;
      write_address_data_log_force[5650] <= 6'h00;
      write_address_data_log_force[5651] <= 6'h00;
      write_address_data_log_force[5652] <= 6'h00;
      write_address_data_log_force[5653] <= 6'h00;
      write_address_data_log_force[5654] <= 6'h00;
      write_address_data_log_force[5655] <= 6'h00;
      write_address_data_log_force[5656] <= 6'h00;
      write_address_data_log_force[5657] <= 6'h00;
      write_address_data_log_force[5658] <= 6'h00;
      write_address_data_log_force[5659] <= 6'h00;
      write_address_data_log_force[5660] <= 6'h00;
      write_address_data_log_force[5661] <= 6'h00;
      write_address_data_log_force[5662] <= 6'h00;
      write_address_data_log_force[5663] <= 6'h00;
      write_address_data_log_force[5664] <= 6'h00;
      write_address_data_log_force[5665] <= 6'h00;
      write_address_data_log_force[5666] <= 6'h00;
      write_address_data_log_force[5667] <= 6'h00;
      write_address_data_log_force[5668] <= 6'h00;
      write_address_data_log_force[5669] <= 6'h00;
      write_address_data_log_force[5670] <= 6'h00;
      write_address_data_log_force[5671] <= 6'h00;
      write_address_data_log_force[5672] <= 6'h00;
      write_address_data_log_force[5673] <= 6'h00;
      write_address_data_log_force[5674] <= 6'h00;
      write_address_data_log_force[5675] <= 6'h00;
      write_address_data_log_force[5676] <= 6'h00;
      write_address_data_log_force[5677] <= 6'h00;
      write_address_data_log_force[5678] <= 6'h00;
      write_address_data_log_force[5679] <= 6'h00;
      write_address_data_log_force[5680] <= 6'h00;
      write_address_data_log_force[5681] <= 6'h00;
      write_address_data_log_force[5682] <= 6'h00;
      write_address_data_log_force[5683] <= 6'h00;
      write_address_data_log_force[5684] <= 6'h00;
      write_address_data_log_force[5685] <= 6'h00;
      write_address_data_log_force[5686] <= 6'h00;
      write_address_data_log_force[5687] <= 6'h00;
      write_address_data_log_force[5688] <= 6'h00;
      write_address_data_log_force[5689] <= 6'h00;
      write_address_data_log_force[5690] <= 6'h00;
      write_address_data_log_force[5691] <= 6'h00;
      write_address_data_log_force[5692] <= 6'h00;
      write_address_data_log_force[5693] <= 6'h00;
      write_address_data_log_force[5694] <= 6'h00;
      write_address_data_log_force[5695] <= 6'h00;
      write_address_data_log_force[5696] <= 6'h00;
      write_address_data_log_force[5697] <= 6'h00;
      write_address_data_log_force[5698] <= 6'h00;
      write_address_data_log_force[5699] <= 6'h00;
      write_address_data_log_force[5700] <= 6'h00;
      write_address_data_log_force[5701] <= 6'h00;
      write_address_data_log_force[5702] <= 6'h00;
      write_address_data_log_force[5703] <= 6'h00;
      write_address_data_log_force[5704] <= 6'h00;
      write_address_data_log_force[5705] <= 6'h00;
      write_address_data_log_force[5706] <= 6'h00;
      write_address_data_log_force[5707] <= 6'h00;
      write_address_data_log_force[5708] <= 6'h00;
      write_address_data_log_force[5709] <= 6'h00;
      write_address_data_log_force[5710] <= 6'h00;
      write_address_data_log_force[5711] <= 6'h00;
      write_address_data_log_force[5712] <= 6'h00;
      write_address_data_log_force[5713] <= 6'h00;
      write_address_data_log_force[5714] <= 6'h00;
      write_address_data_log_force[5715] <= 6'h00;
      write_address_data_log_force[5716] <= 6'h00;
      write_address_data_log_force[5717] <= 6'h00;
      write_address_data_log_force[5718] <= 6'h00;
      write_address_data_log_force[5719] <= 6'h00;
      write_address_data_log_force[5720] <= 6'h00;
      write_address_data_log_force[5721] <= 6'h00;
      write_address_data_log_force[5722] <= 6'h00;
      write_address_data_log_force[5723] <= 6'h00;
      write_address_data_log_force[5724] <= 6'h00;
      write_address_data_log_force[5725] <= 6'h00;
      write_address_data_log_force[5726] <= 6'h00;
      write_address_data_log_force[5727] <= 6'h00;
      write_address_data_log_force[5728] <= 6'h00;
      write_address_data_log_force[5729] <= 6'h00;
      write_address_data_log_force[5730] <= 6'h00;
      write_address_data_log_force[5731] <= 6'h00;
      write_address_data_log_force[5732] <= 6'h00;
      write_address_data_log_force[5733] <= 6'h00;
      write_address_data_log_force[5734] <= 6'h00;
      write_address_data_log_force[5735] <= 6'h00;
      write_address_data_log_force[5736] <= 6'h00;
      write_address_data_log_force[5737] <= 6'h00;
      write_address_data_log_force[5738] <= 6'h00;
      write_address_data_log_force[5739] <= 6'h00;
      write_address_data_log_force[5740] <= 6'h00;
      write_address_data_log_force[5741] <= 6'h00;
      write_address_data_log_force[5742] <= 6'h00;
      write_address_data_log_force[5743] <= 6'h00;
      write_address_data_log_force[5744] <= 6'h00;
      write_address_data_log_force[5745] <= 6'h00;
      write_address_data_log_force[5746] <= 6'h00;
      write_address_data_log_force[5747] <= 6'h00;
      write_address_data_log_force[5748] <= 6'h00;
      write_address_data_log_force[5749] <= 6'h00;
      write_address_data_log_force[5750] <= 6'h00;
      write_address_data_log_force[5751] <= 6'h00;
      write_address_data_log_force[5752] <= 6'h00;
      write_address_data_log_force[5753] <= 6'h00;
      write_address_data_log_force[5754] <= 6'h00;
      write_address_data_log_force[5755] <= 6'h00;
      write_address_data_log_force[5756] <= 6'h00;
      write_address_data_log_force[5757] <= 6'h00;
      write_address_data_log_force[5758] <= 6'h00;
      write_address_data_log_force[5759] <= 6'h00;
      write_address_data_log_force[5760] <= 6'h00;
      write_address_data_log_force[5761] <= 6'h00;
      write_address_data_log_force[5762] <= 6'h00;
      write_address_data_log_force[5763] <= 6'h00;
      write_address_data_log_force[5764] <= 6'h00;
      write_address_data_log_force[5765] <= 6'h00;
      write_address_data_log_force[5766] <= 6'h00;
      write_address_data_log_force[5767] <= 6'h00;
      write_address_data_log_force[5768] <= 6'h00;
      write_address_data_log_force[5769] <= 6'h00;
      write_address_data_log_force[5770] <= 6'h00;
      write_address_data_log_force[5771] <= 6'h00;
      write_address_data_log_force[5772] <= 6'h00;
      write_address_data_log_force[5773] <= 6'h00;
      write_address_data_log_force[5774] <= 6'h00;
      write_address_data_log_force[5775] <= 6'h00;
      write_address_data_log_force[5776] <= 6'h00;
      write_address_data_log_force[5777] <= 6'h00;
      write_address_data_log_force[5778] <= 6'h00;
      write_address_data_log_force[5779] <= 6'h00;
      write_address_data_log_force[5780] <= 6'h00;
      write_address_data_log_force[5781] <= 6'h00;
      write_address_data_log_force[5782] <= 6'h00;
      write_address_data_log_force[5783] <= 6'h00;
      write_address_data_log_force[5784] <= 6'h00;
      write_address_data_log_force[5785] <= 6'h00;
      write_address_data_log_force[5786] <= 6'h00;
      write_address_data_log_force[5787] <= 6'h00;
      write_address_data_log_force[5788] <= 6'h00;
      write_address_data_log_force[5789] <= 6'h00;
      write_address_data_log_force[5790] <= 6'h00;
      write_address_data_log_force[5791] <= 6'h00;
      write_address_data_log_force[5792] <= 6'h00;
      write_address_data_log_force[5793] <= 6'h00;
      write_address_data_log_force[5794] <= 6'h00;
      write_address_data_log_force[5795] <= 6'h00;
      write_address_data_log_force[5796] <= 6'h00;
      write_address_data_log_force[5797] <= 6'h00;
      write_address_data_log_force[5798] <= 6'h00;
      write_address_data_log_force[5799] <= 6'h00;
      write_address_data_log_force[5800] <= 6'h00;
      write_address_data_log_force[5801] <= 6'h00;
      write_address_data_log_force[5802] <= 6'h00;
      write_address_data_log_force[5803] <= 6'h00;
      write_address_data_log_force[5804] <= 6'h00;
      write_address_data_log_force[5805] <= 6'h00;
      write_address_data_log_force[5806] <= 6'h00;
      write_address_data_log_force[5807] <= 6'h00;
      write_address_data_log_force[5808] <= 6'h00;
      write_address_data_log_force[5809] <= 6'h00;
      write_address_data_log_force[5810] <= 6'h00;
      write_address_data_log_force[5811] <= 6'h00;
      write_address_data_log_force[5812] <= 6'h00;
      write_address_data_log_force[5813] <= 6'h00;
      write_address_data_log_force[5814] <= 6'h00;
      write_address_data_log_force[5815] <= 6'h00;
      write_address_data_log_force[5816] <= 6'h00;
      write_address_data_log_force[5817] <= 6'h00;
      write_address_data_log_force[5818] <= 6'h00;
      write_address_data_log_force[5819] <= 6'h00;
      write_address_data_log_force[5820] <= 6'h00;
      write_address_data_log_force[5821] <= 6'h00;
      write_address_data_log_force[5822] <= 6'h00;
      write_address_data_log_force[5823] <= 6'h00;
      write_address_data_log_force[5824] <= 6'h00;
      write_address_data_log_force[5825] <= 6'h00;
      write_address_data_log_force[5826] <= 6'h00;
      write_address_data_log_force[5827] <= 6'h00;
      write_address_data_log_force[5828] <= 6'h00;
      write_address_data_log_force[5829] <= 6'h00;
      write_address_data_log_force[5830] <= 6'h00;
      write_address_data_log_force[5831] <= 6'h00;
      write_address_data_log_force[5832] <= 6'h00;
      write_address_data_log_force[5833] <= 6'h00;
      write_address_data_log_force[5834] <= 6'h00;
      write_address_data_log_force[5835] <= 6'h00;
      write_address_data_log_force[5836] <= 6'h00;
      write_address_data_log_force[5837] <= 6'h00;
      write_address_data_log_force[5838] <= 6'h00;
      write_address_data_log_force[5839] <= 6'h00;
      write_address_data_log_force[5840] <= 6'h00;
      write_address_data_log_force[5841] <= 6'h00;
      write_address_data_log_force[5842] <= 6'h00;
      write_address_data_log_force[5843] <= 6'h00;
      write_address_data_log_force[5844] <= 6'h00;
      write_address_data_log_force[5845] <= 6'h00;
      write_address_data_log_force[5846] <= 6'h00;
      write_address_data_log_force[5847] <= 6'h00;
      write_address_data_log_force[5848] <= 6'h00;
      write_address_data_log_force[5849] <= 6'h00;
      write_address_data_log_force[5850] <= 6'h00;
      write_address_data_log_force[5851] <= 6'h00;
      write_address_data_log_force[5852] <= 6'h00;
      write_address_data_log_force[5853] <= 6'h00;
      write_address_data_log_force[5854] <= 6'h00;
      write_address_data_log_force[5855] <= 6'h00;
      write_address_data_log_force[5856] <= 6'h00;
      write_address_data_log_force[5857] <= 6'h00;
      write_address_data_log_force[5858] <= 6'h00;
      write_address_data_log_force[5859] <= 6'h00;
      write_address_data_log_force[5860] <= 6'h00;
      write_address_data_log_force[5861] <= 6'h00;
      write_address_data_log_force[5862] <= 6'h00;
      write_address_data_log_force[5863] <= 6'h00;
      write_address_data_log_force[5864] <= 6'h00;
      write_address_data_log_force[5865] <= 6'h00;
      write_address_data_log_force[5866] <= 6'h00;
      write_address_data_log_force[5867] <= 6'h00;
      write_address_data_log_force[5868] <= 6'h00;
      write_address_data_log_force[5869] <= 6'h00;
      write_address_data_log_force[5870] <= 6'h00;
      write_address_data_log_force[5871] <= 6'h00;
      write_address_data_log_force[5872] <= 6'h00;
      write_address_data_log_force[5873] <= 6'h00;
      write_address_data_log_force[5874] <= 6'h00;
      write_address_data_log_force[5875] <= 6'h00;
      write_address_data_log_force[5876] <= 6'h00;
      write_address_data_log_force[5877] <= 6'h00;
      write_address_data_log_force[5878] <= 6'h00;
      write_address_data_log_force[5879] <= 6'h00;
      write_address_data_log_force[5880] <= 6'h00;
      write_address_data_log_force[5881] <= 6'h00;
      write_address_data_log_force[5882] <= 6'h00;
      write_address_data_log_force[5883] <= 6'h00;
      write_address_data_log_force[5884] <= 6'h00;
      write_address_data_log_force[5885] <= 6'h00;
      write_address_data_log_force[5886] <= 6'h00;
      write_address_data_log_force[5887] <= 6'h00;
      write_address_data_log_force[5888] <= 6'h00;
      write_address_data_log_force[5889] <= 6'h00;
      write_address_data_log_force[5890] <= 6'h00;
      write_address_data_log_force[5891] <= 6'h00;
      write_address_data_log_force[5892] <= 6'h00;
      write_address_data_log_force[5893] <= 6'h00;
      write_address_data_log_force[5894] <= 6'h00;
      write_address_data_log_force[5895] <= 6'h00;
      write_address_data_log_force[5896] <= 6'h00;
      write_address_data_log_force[5897] <= 6'h00;
      write_address_data_log_force[5898] <= 6'h00;
      write_address_data_log_force[5899] <= 6'h00;
      write_address_data_log_force[5900] <= 6'h00;
      write_address_data_log_force[5901] <= 6'h00;
      write_address_data_log_force[5902] <= 6'h00;
      write_address_data_log_force[5903] <= 6'h00;
      write_address_data_log_force[5904] <= 6'h00;
      write_address_data_log_force[5905] <= 6'h00;
      write_address_data_log_force[5906] <= 6'h00;
      write_address_data_log_force[5907] <= 6'h00;
      write_address_data_log_force[5908] <= 6'h00;
      write_address_data_log_force[5909] <= 6'h00;
      write_address_data_log_force[5910] <= 6'h00;
      write_address_data_log_force[5911] <= 6'h00;
      write_address_data_log_force[5912] <= 6'h00;
      write_address_data_log_force[5913] <= 6'h00;
      write_address_data_log_force[5914] <= 6'h00;
      write_address_data_log_force[5915] <= 6'h00;
      write_address_data_log_force[5916] <= 6'h00;
      write_address_data_log_force[5917] <= 6'h00;
      write_address_data_log_force[5918] <= 6'h00;
      write_address_data_log_force[5919] <= 6'h00;
      write_address_data_log_force[5920] <= 6'h00;
      write_address_data_log_force[5921] <= 6'h00;
      write_address_data_log_force[5922] <= 6'h00;
      write_address_data_log_force[5923] <= 6'h00;
      write_address_data_log_force[5924] <= 6'h00;
      write_address_data_log_force[5925] <= 6'h00;
      write_address_data_log_force[5926] <= 6'h00;
      write_address_data_log_force[5927] <= 6'h00;
      write_address_data_log_force[5928] <= 6'h00;
      write_address_data_log_force[5929] <= 6'h00;
      write_address_data_log_force[5930] <= 6'h00;
      write_address_data_log_force[5931] <= 6'h00;
      write_address_data_log_force[5932] <= 6'h00;
      write_address_data_log_force[5933] <= 6'h00;
      write_address_data_log_force[5934] <= 6'h00;
      write_address_data_log_force[5935] <= 6'h00;
      write_address_data_log_force[5936] <= 6'h00;
      write_address_data_log_force[5937] <= 6'h00;
      write_address_data_log_force[5938] <= 6'h00;
      write_address_data_log_force[5939] <= 6'h00;
      write_address_data_log_force[5940] <= 6'h00;
      write_address_data_log_force[5941] <= 6'h00;
      write_address_data_log_force[5942] <= 6'h00;
      write_address_data_log_force[5943] <= 6'h00;
      write_address_data_log_force[5944] <= 6'h00;
      write_address_data_log_force[5945] <= 6'h00;
      write_address_data_log_force[5946] <= 6'h00;
      write_address_data_log_force[5947] <= 6'h00;
      write_address_data_log_force[5948] <= 6'h00;
      write_address_data_log_force[5949] <= 6'h00;
      write_address_data_log_force[5950] <= 6'h00;
      write_address_data_log_force[5951] <= 6'h00;
      write_address_data_log_force[5952] <= 6'h00;
      write_address_data_log_force[5953] <= 6'h00;
      write_address_data_log_force[5954] <= 6'h00;
      write_address_data_log_force[5955] <= 6'h00;
      write_address_data_log_force[5956] <= 6'h00;
      write_address_data_log_force[5957] <= 6'h00;
      write_address_data_log_force[5958] <= 6'h00;
      write_address_data_log_force[5959] <= 6'h00;
      write_address_data_log_force[5960] <= 6'h00;
      write_address_data_log_force[5961] <= 6'h00;
      write_address_data_log_force[5962] <= 6'h00;
      write_address_data_log_force[5963] <= 6'h00;
      write_address_data_log_force[5964] <= 6'h00;
      write_address_data_log_force[5965] <= 6'h00;
      write_address_data_log_force[5966] <= 6'h00;
      write_address_data_log_force[5967] <= 6'h00;
      write_address_data_log_force[5968] <= 6'h00;
      write_address_data_log_force[5969] <= 6'h00;
      write_address_data_log_force[5970] <= 6'h00;
      write_address_data_log_force[5971] <= 6'h00;
      write_address_data_log_force[5972] <= 6'h00;
      write_address_data_log_force[5973] <= 6'h00;
      write_address_data_log_force[5974] <= 6'h00;
      write_address_data_log_force[5975] <= 6'h00;
      write_address_data_log_force[5976] <= 6'h00;
      write_address_data_log_force[5977] <= 6'h00;
      write_address_data_log_force[5978] <= 6'h00;
      write_address_data_log_force[5979] <= 6'h00;
      write_address_data_log_force[5980] <= 6'h00;
      write_address_data_log_force[5981] <= 6'h00;
      write_address_data_log_force[5982] <= 6'h00;
      write_address_data_log_force[5983] <= 6'h00;
      write_address_data_log_force[5984] <= 6'h00;
      write_address_data_log_force[5985] <= 6'h00;
      write_address_data_log_force[5986] <= 6'h00;
      write_address_data_log_force[5987] <= 6'h00;
      write_address_data_log_force[5988] <= 6'h00;
      write_address_data_log_force[5989] <= 6'h00;
      write_address_data_log_force[5990] <= 6'h00;
      write_address_data_log_force[5991] <= 6'h00;
      write_address_data_log_force[5992] <= 6'h00;
      write_address_data_log_force[5993] <= 6'h00;
      write_address_data_log_force[5994] <= 6'h00;
      write_address_data_log_force[5995] <= 6'h00;
      write_address_data_log_force[5996] <= 6'h00;
      write_address_data_log_force[5997] <= 6'h00;
      write_address_data_log_force[5998] <= 6'h00;
      write_address_data_log_force[5999] <= 6'h00;
      write_address_data_log_force[6000] <= 6'h00;
      write_address_data_log_force[6001] <= 6'h00;
      write_address_data_log_force[6002] <= 6'h00;
      write_address_data_log_force[6003] <= 6'h00;
      write_address_data_log_force[6004] <= 6'h00;
      write_address_data_log_force[6005] <= 6'h00;
      write_address_data_log_force[6006] <= 6'h00;
      write_address_data_log_force[6007] <= 6'h00;
      write_address_data_log_force[6008] <= 6'h00;
      write_address_data_log_force[6009] <= 6'h00;
      write_address_data_log_force[6010] <= 6'h00;
      write_address_data_log_force[6011] <= 6'h00;
      write_address_data_log_force[6012] <= 6'h00;
      write_address_data_log_force[6013] <= 6'h00;
      write_address_data_log_force[6014] <= 6'h00;
      write_address_data_log_force[6015] <= 6'h00;
      write_address_data_log_force[6016] <= 6'h00;
      write_address_data_log_force[6017] <= 6'h00;
      write_address_data_log_force[6018] <= 6'h00;
      write_address_data_log_force[6019] <= 6'h00;
      write_address_data_log_force[6020] <= 6'h00;
      write_address_data_log_force[6021] <= 6'h00;
      write_address_data_log_force[6022] <= 6'h00;
      write_address_data_log_force[6023] <= 6'h00;
      write_address_data_log_force[6024] <= 6'h00;
      write_address_data_log_force[6025] <= 6'h00;
      write_address_data_log_force[6026] <= 6'h00;
      write_address_data_log_force[6027] <= 6'h00;
      write_address_data_log_force[6028] <= 6'h00;
      write_address_data_log_force[6029] <= 6'h00;
      write_address_data_log_force[6030] <= 6'h00;
      write_address_data_log_force[6031] <= 6'h00;
      write_address_data_log_force[6032] <= 6'h00;
      write_address_data_log_force[6033] <= 6'h00;
      write_address_data_log_force[6034] <= 6'h00;
      write_address_data_log_force[6035] <= 6'h00;
      write_address_data_log_force[6036] <= 6'h00;
      write_address_data_log_force[6037] <= 6'h00;
      write_address_data_log_force[6038] <= 6'h00;
      write_address_data_log_force[6039] <= 6'h00;
      write_address_data_log_force[6040] <= 6'h00;
      write_address_data_log_force[6041] <= 6'h00;
      write_address_data_log_force[6042] <= 6'h00;
      write_address_data_log_force[6043] <= 6'h00;
      write_address_data_log_force[6044] <= 6'h00;
      write_address_data_log_force[6045] <= 6'h00;
      write_address_data_log_force[6046] <= 6'h00;
      write_address_data_log_force[6047] <= 6'h00;
      write_address_data_log_force[6048] <= 6'h00;
      write_address_data_log_force[6049] <= 6'h00;
      write_address_data_log_force[6050] <= 6'h00;
      write_address_data_log_force[6051] <= 6'h00;
      write_address_data_log_force[6052] <= 6'h00;
      write_address_data_log_force[6053] <= 6'h00;
      write_address_data_log_force[6054] <= 6'h00;
      write_address_data_log_force[6055] <= 6'h00;
      write_address_data_log_force[6056] <= 6'h00;
      write_address_data_log_force[6057] <= 6'h00;
      write_address_data_log_force[6058] <= 6'h00;
      write_address_data_log_force[6059] <= 6'h00;
      write_address_data_log_force[6060] <= 6'h00;
      write_address_data_log_force[6061] <= 6'h00;
      write_address_data_log_force[6062] <= 6'h00;
      write_address_data_log_force[6063] <= 6'h00;
      write_address_data_log_force[6064] <= 6'h00;
      write_address_data_log_force[6065] <= 6'h00;
      write_address_data_log_force[6066] <= 6'h00;
      write_address_data_log_force[6067] <= 6'h00;
      write_address_data_log_force[6068] <= 6'h00;
      write_address_data_log_force[6069] <= 6'h00;
      write_address_data_log_force[6070] <= 6'h00;
      write_address_data_log_force[6071] <= 6'h00;
      write_address_data_log_force[6072] <= 6'h00;
      write_address_data_log_force[6073] <= 6'h00;
      write_address_data_log_force[6074] <= 6'h00;
      write_address_data_log_force[6075] <= 6'h00;
      write_address_data_log_force[6076] <= 6'h00;
      write_address_data_log_force[6077] <= 6'h00;
      write_address_data_log_force[6078] <= 6'h00;
      write_address_data_log_force[6079] <= 6'h00;
      write_address_data_log_force[6080] <= 6'h00;
      write_address_data_log_force[6081] <= 6'h00;
      write_address_data_log_force[6082] <= 6'h00;
      write_address_data_log_force[6083] <= 6'h00;
      write_address_data_log_force[6084] <= 6'h00;
      write_address_data_log_force[6085] <= 6'h00;
      write_address_data_log_force[6086] <= 6'h00;
      write_address_data_log_force[6087] <= 6'h00;
      write_address_data_log_force[6088] <= 6'h00;
      write_address_data_log_force[6089] <= 6'h00;
      write_address_data_log_force[6090] <= 6'h00;
      write_address_data_log_force[6091] <= 6'h00;
      write_address_data_log_force[6092] <= 6'h00;
      write_address_data_log_force[6093] <= 6'h00;
      write_address_data_log_force[6094] <= 6'h00;
      write_address_data_log_force[6095] <= 6'h00;
      write_address_data_log_force[6096] <= 6'h00;
      write_address_data_log_force[6097] <= 6'h00;
      write_address_data_log_force[6098] <= 6'h00;
      write_address_data_log_force[6099] <= 6'h00;
      write_address_data_log_force[6100] <= 6'h00;
      write_address_data_log_force[6101] <= 6'h00;
      write_address_data_log_force[6102] <= 6'h00;
      write_address_data_log_force[6103] <= 6'h00;
      write_address_data_log_force[6104] <= 6'h00;
      write_address_data_log_force[6105] <= 6'h00;
      write_address_data_log_force[6106] <= 6'h00;
      write_address_data_log_force[6107] <= 6'h00;
      write_address_data_log_force[6108] <= 6'h00;
      write_address_data_log_force[6109] <= 6'h00;
      write_address_data_log_force[6110] <= 6'h00;
      write_address_data_log_force[6111] <= 6'h00;
      write_address_data_log_force[6112] <= 6'h00;
      write_address_data_log_force[6113] <= 6'h00;
      write_address_data_log_force[6114] <= 6'h00;
      write_address_data_log_force[6115] <= 6'h00;
      write_address_data_log_force[6116] <= 6'h00;
      write_address_data_log_force[6117] <= 6'h00;
      write_address_data_log_force[6118] <= 6'h00;
      write_address_data_log_force[6119] <= 6'h00;
      write_address_data_log_force[6120] <= 6'h00;
      write_address_data_log_force[6121] <= 6'h00;
      write_address_data_log_force[6122] <= 6'h00;
      write_address_data_log_force[6123] <= 6'h00;
      write_address_data_log_force[6124] <= 6'h00;
      write_address_data_log_force[6125] <= 6'h00;
      write_address_data_log_force[6126] <= 6'h00;
      write_address_data_log_force[6127] <= 6'h00;
      write_address_data_log_force[6128] <= 6'h00;
      write_address_data_log_force[6129] <= 6'h00;
      write_address_data_log_force[6130] <= 6'h00;
      write_address_data_log_force[6131] <= 6'h00;
      write_address_data_log_force[6132] <= 6'h00;
      write_address_data_log_force[6133] <= 6'h00;
      write_address_data_log_force[6134] <= 6'h00;
      write_address_data_log_force[6135] <= 6'h00;
      write_address_data_log_force[6136] <= 6'h00;
      write_address_data_log_force[6137] <= 6'h00;
      write_address_data_log_force[6138] <= 6'h00;
      write_address_data_log_force[6139] <= 6'h00;
      write_address_data_log_force[6140] <= 6'h00;
      write_address_data_log_force[6141] <= 6'h00;
      write_address_data_log_force[6142] <= 6'h00;
      write_address_data_log_force[6143] <= 6'h00;
      write_address_data_log_force[6144] <= 6'h00;
      write_address_data_log_force[6145] <= 6'h00;
      write_address_data_log_force[6146] <= 6'h00;
      write_address_data_log_force[6147] <= 6'h00;
      write_address_data_log_force[6148] <= 6'h00;
      write_address_data_log_force[6149] <= 6'h00;
      write_address_data_log_force[6150] <= 6'h00;
      write_address_data_log_force[6151] <= 6'h00;
      write_address_data_log_force[6152] <= 6'h00;
      write_address_data_log_force[6153] <= 6'h00;
      write_address_data_log_force[6154] <= 6'h00;
      write_address_data_log_force[6155] <= 6'h00;
      write_address_data_log_force[6156] <= 6'h00;
      write_address_data_log_force[6157] <= 6'h00;
      write_address_data_log_force[6158] <= 6'h00;
      write_address_data_log_force[6159] <= 6'h00;
      write_address_data_log_force[6160] <= 6'h00;
      write_address_data_log_force[6161] <= 6'h00;
      write_address_data_log_force[6162] <= 6'h00;
      write_address_data_log_force[6163] <= 6'h00;
      write_address_data_log_force[6164] <= 6'h00;
      write_address_data_log_force[6165] <= 6'h00;
      write_address_data_log_force[6166] <= 6'h00;
      write_address_data_log_force[6167] <= 6'h00;
      write_address_data_log_force[6168] <= 6'h00;
      write_address_data_log_force[6169] <= 6'h00;
      write_address_data_log_force[6170] <= 6'h00;
      write_address_data_log_force[6171] <= 6'h00;
      write_address_data_log_force[6172] <= 6'h00;
      write_address_data_log_force[6173] <= 6'h00;
      write_address_data_log_force[6174] <= 6'h00;
      write_address_data_log_force[6175] <= 6'h00;
      write_address_data_log_force[6176] <= 6'h00;
      write_address_data_log_force[6177] <= 6'h00;
      write_address_data_log_force[6178] <= 6'h00;
      write_address_data_log_force[6179] <= 6'h00;
      write_address_data_log_force[6180] <= 6'h00;
      write_address_data_log_force[6181] <= 6'h00;
      write_address_data_log_force[6182] <= 6'h00;
      write_address_data_log_force[6183] <= 6'h00;
      write_address_data_log_force[6184] <= 6'h00;
      write_address_data_log_force[6185] <= 6'h00;
      write_address_data_log_force[6186] <= 6'h00;
      write_address_data_log_force[6187] <= 6'h00;
      write_address_data_log_force[6188] <= 6'h00;
      write_address_data_log_force[6189] <= 6'h00;
      write_address_data_log_force[6190] <= 6'h00;
      write_address_data_log_force[6191] <= 6'h00;
      write_address_data_log_force[6192] <= 6'h00;
      write_address_data_log_force[6193] <= 6'h00;
      write_address_data_log_force[6194] <= 6'h00;
      write_address_data_log_force[6195] <= 6'h00;
      write_address_data_log_force[6196] <= 6'h00;
      write_address_data_log_force[6197] <= 6'h00;
      write_address_data_log_force[6198] <= 6'h00;
      write_address_data_log_force[6199] <= 6'h00;
      write_address_data_log_force[6200] <= 6'h00;
      write_address_data_log_force[6201] <= 6'h00;
      write_address_data_log_force[6202] <= 6'h00;
      write_address_data_log_force[6203] <= 6'h00;
      write_address_data_log_force[6204] <= 6'h00;
      write_address_data_log_force[6205] <= 6'h00;
      write_address_data_log_force[6206] <= 6'h00;
      write_address_data_log_force[6207] <= 6'h00;
      write_address_data_log_force[6208] <= 6'h00;
      write_address_data_log_force[6209] <= 6'h00;
      write_address_data_log_force[6210] <= 6'h00;
      write_address_data_log_force[6211] <= 6'h00;
      write_address_data_log_force[6212] <= 6'h00;
      write_address_data_log_force[6213] <= 6'h00;
      write_address_data_log_force[6214] <= 6'h00;
      write_address_data_log_force[6215] <= 6'h00;
      write_address_data_log_force[6216] <= 6'h00;
      write_address_data_log_force[6217] <= 6'h00;
      write_address_data_log_force[6218] <= 6'h00;
      write_address_data_log_force[6219] <= 6'h00;
      write_address_data_log_force[6220] <= 6'h00;
      write_address_data_log_force[6221] <= 6'h00;
      write_address_data_log_force[6222] <= 6'h00;
      write_address_data_log_force[6223] <= 6'h00;
      write_address_data_log_force[6224] <= 6'h00;
      write_address_data_log_force[6225] <= 6'h00;
      write_address_data_log_force[6226] <= 6'h00;
      write_address_data_log_force[6227] <= 6'h00;
      write_address_data_log_force[6228] <= 6'h00;
      write_address_data_log_force[6229] <= 6'h00;
      write_address_data_log_force[6230] <= 6'h00;
      write_address_data_log_force[6231] <= 6'h00;
      write_address_data_log_force[6232] <= 6'h00;
      write_address_data_log_force[6233] <= 6'h00;
      write_address_data_log_force[6234] <= 6'h00;
      write_address_data_log_force[6235] <= 6'h00;
      write_address_data_log_force[6236] <= 6'h00;
      write_address_data_log_force[6237] <= 6'h00;
      write_address_data_log_force[6238] <= 6'h00;
      write_address_data_log_force[6239] <= 6'h00;
      write_address_data_log_force[6240] <= 6'h00;
      write_address_data_log_force[6241] <= 6'h00;
      write_address_data_log_force[6242] <= 6'h00;
      write_address_data_log_force[6243] <= 6'h00;
      write_address_data_log_force[6244] <= 6'h00;
      write_address_data_log_force[6245] <= 6'h00;
      write_address_data_log_force[6246] <= 6'h00;
      write_address_data_log_force[6247] <= 6'h00;
      write_address_data_log_force[6248] <= 6'h00;
      write_address_data_log_force[6249] <= 6'h00;
      write_address_data_log_force[6250] <= 6'h00;
      write_address_data_log_force[6251] <= 6'h00;
      write_address_data_log_force[6252] <= 6'h00;
      write_address_data_log_force[6253] <= 6'h00;
      write_address_data_log_force[6254] <= 6'h00;
      write_address_data_log_force[6255] <= 6'h00;
      write_address_data_log_force[6256] <= 6'h00;
      write_address_data_log_force[6257] <= 6'h00;
      write_address_data_log_force[6258] <= 6'h00;
      write_address_data_log_force[6259] <= 6'h00;
      write_address_data_log_force[6260] <= 6'h00;
      write_address_data_log_force[6261] <= 6'h00;
      write_address_data_log_force[6262] <= 6'h00;
      write_address_data_log_force[6263] <= 6'h00;
      write_address_data_log_force[6264] <= 6'h00;
      write_address_data_log_force[6265] <= 6'h00;
      write_address_data_log_force[6266] <= 6'h00;
      write_address_data_log_force[6267] <= 6'h00;
      write_address_data_log_force[6268] <= 6'h00;
      write_address_data_log_force[6269] <= 6'h00;
      write_address_data_log_force[6270] <= 6'h00;
      write_address_data_log_force[6271] <= 6'h00;
      write_address_data_log_force[6272] <= 6'h00;
      write_address_data_log_force[6273] <= 6'h00;
      write_address_data_log_force[6274] <= 6'h00;
      write_address_data_log_force[6275] <= 6'h00;
      write_address_data_log_force[6276] <= 6'h00;
      write_address_data_log_force[6277] <= 6'h00;
      write_address_data_log_force[6278] <= 6'h00;
      write_address_data_log_force[6279] <= 6'h00;
      write_address_data_log_force[6280] <= 6'h00;
      write_address_data_log_force[6281] <= 6'h00;
      write_address_data_log_force[6282] <= 6'h00;
      write_address_data_log_force[6283] <= 6'h00;
      write_address_data_log_force[6284] <= 6'h00;
      write_address_data_log_force[6285] <= 6'h00;
      write_address_data_log_force[6286] <= 6'h00;
      write_address_data_log_force[6287] <= 6'h00;
      write_address_data_log_force[6288] <= 6'h00;
      write_address_data_log_force[6289] <= 6'h00;
      write_address_data_log_force[6290] <= 6'h00;
      write_address_data_log_force[6291] <= 6'h00;
      write_address_data_log_force[6292] <= 6'h00;
      write_address_data_log_force[6293] <= 6'h00;
      write_address_data_log_force[6294] <= 6'h00;
      write_address_data_log_force[6295] <= 6'h00;
      write_address_data_log_force[6296] <= 6'h00;
      write_address_data_log_force[6297] <= 6'h00;
      write_address_data_log_force[6298] <= 6'h00;
      write_address_data_log_force[6299] <= 6'h00;
      write_address_data_log_force[6300] <= 6'h00;
      write_address_data_log_force[6301] <= 6'h00;
      write_address_data_log_force[6302] <= 6'h00;
      write_address_data_log_force[6303] <= 6'h00;
      write_address_data_log_force[6304] <= 6'h00;
      write_address_data_log_force[6305] <= 6'h00;
      write_address_data_log_force[6306] <= 6'h00;
      write_address_data_log_force[6307] <= 6'h00;
      write_address_data_log_force[6308] <= 6'h00;
      write_address_data_log_force[6309] <= 6'h00;
      write_address_data_log_force[6310] <= 6'h00;
      write_address_data_log_force[6311] <= 6'h00;
      write_address_data_log_force[6312] <= 6'h00;
      write_address_data_log_force[6313] <= 6'h00;
      write_address_data_log_force[6314] <= 6'h00;
      write_address_data_log_force[6315] <= 6'h00;
      write_address_data_log_force[6316] <= 6'h00;
      write_address_data_log_force[6317] <= 6'h00;
      write_address_data_log_force[6318] <= 6'h00;
      write_address_data_log_force[6319] <= 6'h00;
      write_address_data_log_force[6320] <= 6'h00;
      write_address_data_log_force[6321] <= 6'h00;
      write_address_data_log_force[6322] <= 6'h00;
      write_address_data_log_force[6323] <= 6'h00;
      write_address_data_log_force[6324] <= 6'h00;
      write_address_data_log_force[6325] <= 6'h00;
      write_address_data_log_force[6326] <= 6'h00;
      write_address_data_log_force[6327] <= 6'h00;
      write_address_data_log_force[6328] <= 6'h00;
      write_address_data_log_force[6329] <= 6'h00;
      write_address_data_log_force[6330] <= 6'h00;
      write_address_data_log_force[6331] <= 6'h00;
      write_address_data_log_force[6332] <= 6'h00;
      write_address_data_log_force[6333] <= 6'h00;
      write_address_data_log_force[6334] <= 6'h00;
      write_address_data_log_force[6335] <= 6'h00;
      write_address_data_log_force[6336] <= 6'h00;
      write_address_data_log_force[6337] <= 6'h00;
      write_address_data_log_force[6338] <= 6'h00;
      write_address_data_log_force[6339] <= 6'h00;
      write_address_data_log_force[6340] <= 6'h00;
      write_address_data_log_force[6341] <= 6'h00;
      write_address_data_log_force[6342] <= 6'h00;
      write_address_data_log_force[6343] <= 6'h00;
      write_address_data_log_force[6344] <= 6'h00;
      write_address_data_log_force[6345] <= 6'h00;
      write_address_data_log_force[6346] <= 6'h00;
      write_address_data_log_force[6347] <= 6'h00;
      write_address_data_log_force[6348] <= 6'h00;
      write_address_data_log_force[6349] <= 6'h00;
      write_address_data_log_force[6350] <= 6'h00;
      write_address_data_log_force[6351] <= 6'h00;
      write_address_data_log_force[6352] <= 6'h00;
      write_address_data_log_force[6353] <= 6'h00;
      write_address_data_log_force[6354] <= 6'h00;
      write_address_data_log_force[6355] <= 6'h00;
      write_address_data_log_force[6356] <= 6'h00;
      write_address_data_log_force[6357] <= 6'h00;
      write_address_data_log_force[6358] <= 6'h00;
      write_address_data_log_force[6359] <= 6'h00;
      write_address_data_log_force[6360] <= 6'h00;
      write_address_data_log_force[6361] <= 6'h00;
      write_address_data_log_force[6362] <= 6'h00;
      write_address_data_log_force[6363] <= 6'h00;
      write_address_data_log_force[6364] <= 6'h00;
      write_address_data_log_force[6365] <= 6'h00;
      write_address_data_log_force[6366] <= 6'h00;
      write_address_data_log_force[6367] <= 6'h00;
      write_address_data_log_force[6368] <= 6'h00;
      write_address_data_log_force[6369] <= 6'h00;
      write_address_data_log_force[6370] <= 6'h00;
      write_address_data_log_force[6371] <= 6'h00;
      write_address_data_log_force[6372] <= 6'h00;
      write_address_data_log_force[6373] <= 6'h00;
      write_address_data_log_force[6374] <= 6'h00;
      write_address_data_log_force[6375] <= 6'h00;
      write_address_data_log_force[6376] <= 6'h00;
      write_address_data_log_force[6377] <= 6'h00;
      write_address_data_log_force[6378] <= 6'h00;
      write_address_data_log_force[6379] <= 6'h00;
      write_address_data_log_force[6380] <= 6'h00;
      write_address_data_log_force[6381] <= 6'h00;
      write_address_data_log_force[6382] <= 6'h00;
      write_address_data_log_force[6383] <= 6'h00;
      write_address_data_log_force[6384] <= 6'h00;
      write_address_data_log_force[6385] <= 6'h00;
      write_address_data_log_force[6386] <= 6'h00;
      write_address_data_log_force[6387] <= 6'h00;
      write_address_data_log_force[6388] <= 6'h00;
      write_address_data_log_force[6389] <= 6'h00;
      write_address_data_log_force[6390] <= 6'h00;
      write_address_data_log_force[6391] <= 6'h00;
      write_address_data_log_force[6392] <= 6'h00;
      write_address_data_log_force[6393] <= 6'h00;
      write_address_data_log_force[6394] <= 6'h00;
      write_address_data_log_force[6395] <= 6'h00;
      write_address_data_log_force[6396] <= 6'h00;
      write_address_data_log_force[6397] <= 6'h00;
      write_address_data_log_force[6398] <= 6'h00;
      write_address_data_log_force[6399] <= 6'h00;
      write_address_data_log_force[6400] <= 6'h00;
      write_address_data_log_force[6401] <= 6'h00;
      write_address_data_log_force[6402] <= 6'h00;
      write_address_data_log_force[6403] <= 6'h00;
      write_address_data_log_force[6404] <= 6'h00;
      write_address_data_log_force[6405] <= 6'h00;
      write_address_data_log_force[6406] <= 6'h00;
      write_address_data_log_force[6407] <= 6'h00;
      write_address_data_log_force[6408] <= 6'h00;
      write_address_data_log_force[6409] <= 6'h00;
      write_address_data_log_force[6410] <= 6'h00;
      write_address_data_log_force[6411] <= 6'h00;
      write_address_data_log_force[6412] <= 6'h00;
      write_address_data_log_force[6413] <= 6'h00;
      write_address_data_log_force[6414] <= 6'h00;
      write_address_data_log_force[6415] <= 6'h00;
      write_address_data_log_force[6416] <= 6'h00;
      write_address_data_log_force[6417] <= 6'h00;
      write_address_data_log_force[6418] <= 6'h00;
      write_address_data_log_force[6419] <= 6'h00;
      write_address_data_log_force[6420] <= 6'h00;
      write_address_data_log_force[6421] <= 6'h00;
      write_address_data_log_force[6422] <= 6'h00;
      write_address_data_log_force[6423] <= 6'h00;
      write_address_data_log_force[6424] <= 6'h00;
      write_address_data_log_force[6425] <= 6'h00;
      write_address_data_log_force[6426] <= 6'h00;
      write_address_data_log_force[6427] <= 6'h00;
      write_address_data_log_force[6428] <= 6'h00;
      write_address_data_log_force[6429] <= 6'h00;
      write_address_data_log_force[6430] <= 6'h00;
      write_address_data_log_force[6431] <= 6'h00;
      write_address_data_log_force[6432] <= 6'h00;
      write_address_data_log_force[6433] <= 6'h00;
      write_address_data_log_force[6434] <= 6'h00;
      write_address_data_log_force[6435] <= 6'h00;
      write_address_data_log_force[6436] <= 6'h00;
      write_address_data_log_force[6437] <= 6'h00;
      write_address_data_log_force[6438] <= 6'h00;
      write_address_data_log_force[6439] <= 6'h00;
      write_address_data_log_force[6440] <= 6'h00;
      write_address_data_log_force[6441] <= 6'h00;
      write_address_data_log_force[6442] <= 6'h00;
      write_address_data_log_force[6443] <= 6'h00;
      write_address_data_log_force[6444] <= 6'h00;
      write_address_data_log_force[6445] <= 6'h00;
      write_address_data_log_force[6446] <= 6'h00;
      write_address_data_log_force[6447] <= 6'h00;
      write_address_data_log_force[6448] <= 6'h00;
      write_address_data_log_force[6449] <= 6'h00;
      write_address_data_log_force[6450] <= 6'h00;
      write_address_data_log_force[6451] <= 6'h00;
      write_address_data_log_force[6452] <= 6'h00;
      write_address_data_log_force[6453] <= 6'h00;
      write_address_data_log_force[6454] <= 6'h00;
      write_address_data_log_force[6455] <= 6'h00;
      write_address_data_log_force[6456] <= 6'h00;
      write_address_data_log_force[6457] <= 6'h00;
      write_address_data_log_force[6458] <= 6'h00;
      write_address_data_log_force[6459] <= 6'h00;
      write_address_data_log_force[6460] <= 6'h00;
      write_address_data_log_force[6461] <= 6'h00;
      write_address_data_log_force[6462] <= 6'h00;
      write_address_data_log_force[6463] <= 6'h00;
      write_address_data_log_force[6464] <= 6'h00;
      write_address_data_log_force[6465] <= 6'h00;
      write_address_data_log_force[6466] <= 6'h00;
      write_address_data_log_force[6467] <= 6'h00;
      write_address_data_log_force[6468] <= 6'h00;
      write_address_data_log_force[6469] <= 6'h00;
      write_address_data_log_force[6470] <= 6'h00;
      write_address_data_log_force[6471] <= 6'h00;
      write_address_data_log_force[6472] <= 6'h00;
      write_address_data_log_force[6473] <= 6'h00;
      write_address_data_log_force[6474] <= 6'h00;
      write_address_data_log_force[6475] <= 6'h00;
      write_address_data_log_force[6476] <= 6'h00;
      write_address_data_log_force[6477] <= 6'h00;
      write_address_data_log_force[6478] <= 6'h00;
      write_address_data_log_force[6479] <= 6'h00;
      write_address_data_log_force[6480] <= 6'h00;
      write_address_data_log_force[6481] <= 6'h00;
      write_address_data_log_force[6482] <= 6'h00;
      write_address_data_log_force[6483] <= 6'h00;
      write_address_data_log_force[6484] <= 6'h00;
      write_address_data_log_force[6485] <= 6'h00;
      write_address_data_log_force[6486] <= 6'h00;
      write_address_data_log_force[6487] <= 6'h00;
      write_address_data_log_force[6488] <= 6'h00;
      write_address_data_log_force[6489] <= 6'h00;
      write_address_data_log_force[6490] <= 6'h00;
      write_address_data_log_force[6491] <= 6'h00;
      write_address_data_log_force[6492] <= 6'h00;
      write_address_data_log_force[6493] <= 6'h00;
      write_address_data_log_force[6494] <= 6'h00;
      write_address_data_log_force[6495] <= 6'h00;
      write_address_data_log_force[6496] <= 6'h00;
      write_address_data_log_force[6497] <= 6'h00;
      write_address_data_log_force[6498] <= 6'h00;
      write_address_data_log_force[6499] <= 6'h00;
      write_address_data_log_force[6500] <= 6'h00;
      write_address_data_log_force[6501] <= 6'h00;
      write_address_data_log_force[6502] <= 6'h00;
      write_address_data_log_force[6503] <= 6'h00;
      write_address_data_log_force[6504] <= 6'h00;
      write_address_data_log_force[6505] <= 6'h00;
      write_address_data_log_force[6506] <= 6'h00;
      write_address_data_log_force[6507] <= 6'h00;
      write_address_data_log_force[6508] <= 6'h00;
      write_address_data_log_force[6509] <= 6'h00;
      write_address_data_log_force[6510] <= 6'h00;
      write_address_data_log_force[6511] <= 6'h00;
      write_address_data_log_force[6512] <= 6'h00;
      write_address_data_log_force[6513] <= 6'h00;
      write_address_data_log_force[6514] <= 6'h00;
      write_address_data_log_force[6515] <= 6'h00;
      write_address_data_log_force[6516] <= 6'h00;
      write_address_data_log_force[6517] <= 6'h00;
      write_address_data_log_force[6518] <= 6'h00;
      write_address_data_log_force[6519] <= 6'h00;
      write_address_data_log_force[6520] <= 6'h00;
      write_address_data_log_force[6521] <= 6'h00;
      write_address_data_log_force[6522] <= 6'h00;
      write_address_data_log_force[6523] <= 6'h00;
      write_address_data_log_force[6524] <= 6'h00;
      write_address_data_log_force[6525] <= 6'h00;
      write_address_data_log_force[6526] <= 6'h00;
      write_address_data_log_force[6527] <= 6'h00;
      write_address_data_log_force[6528] <= 6'h00;
      write_address_data_log_force[6529] <= 6'h00;
      write_address_data_log_force[6530] <= 6'h00;
      write_address_data_log_force[6531] <= 6'h00;
      write_address_data_log_force[6532] <= 6'h00;
      write_address_data_log_force[6533] <= 6'h00;
      write_address_data_log_force[6534] <= 6'h00;
      write_address_data_log_force[6535] <= 6'h00;
      write_address_data_log_force[6536] <= 6'h00;
      write_address_data_log_force[6537] <= 6'h00;
      write_address_data_log_force[6538] <= 6'h00;
      write_address_data_log_force[6539] <= 6'h00;
      write_address_data_log_force[6540] <= 6'h00;
      write_address_data_log_force[6541] <= 6'h00;
      write_address_data_log_force[6542] <= 6'h00;
      write_address_data_log_force[6543] <= 6'h00;
      write_address_data_log_force[6544] <= 6'h00;
      write_address_data_log_force[6545] <= 6'h00;
      write_address_data_log_force[6546] <= 6'h00;
      write_address_data_log_force[6547] <= 6'h00;
      write_address_data_log_force[6548] <= 6'h00;
      write_address_data_log_force[6549] <= 6'h00;
      write_address_data_log_force[6550] <= 6'h00;
      write_address_data_log_force[6551] <= 6'h00;
      write_address_data_log_force[6552] <= 6'h00;
      write_address_data_log_force[6553] <= 6'h00;
      write_address_data_log_force[6554] <= 6'h00;
      write_address_data_log_force[6555] <= 6'h00;
      write_address_data_log_force[6556] <= 6'h00;
      write_address_data_log_force[6557] <= 6'h00;
      write_address_data_log_force[6558] <= 6'h00;
      write_address_data_log_force[6559] <= 6'h00;
      write_address_data_log_force[6560] <= 6'h00;
      write_address_data_log_force[6561] <= 6'h00;
      write_address_data_log_force[6562] <= 6'h00;
      write_address_data_log_force[6563] <= 6'h00;
      write_address_data_log_force[6564] <= 6'h00;
      write_address_data_log_force[6565] <= 6'h00;
      write_address_data_log_force[6566] <= 6'h00;
      write_address_data_log_force[6567] <= 6'h00;
      write_address_data_log_force[6568] <= 6'h00;
      write_address_data_log_force[6569] <= 6'h00;
      write_address_data_log_force[6570] <= 6'h00;
      write_address_data_log_force[6571] <= 6'h00;
      write_address_data_log_force[6572] <= 6'h00;
      write_address_data_log_force[6573] <= 6'h00;
      write_address_data_log_force[6574] <= 6'h00;
      write_address_data_log_force[6575] <= 6'h00;
      write_address_data_log_force[6576] <= 6'h00;
      write_address_data_log_force[6577] <= 6'h00;
      write_address_data_log_force[6578] <= 6'h00;
      write_address_data_log_force[6579] <= 6'h00;
      write_address_data_log_force[6580] <= 6'h00;
      write_address_data_log_force[6581] <= 6'h00;
      write_address_data_log_force[6582] <= 6'h00;
      write_address_data_log_force[6583] <= 6'h00;
      write_address_data_log_force[6584] <= 6'h00;
      write_address_data_log_force[6585] <= 6'h00;
      write_address_data_log_force[6586] <= 6'h00;
      write_address_data_log_force[6587] <= 6'h00;
      write_address_data_log_force[6588] <= 6'h00;
      write_address_data_log_force[6589] <= 6'h00;
      write_address_data_log_force[6590] <= 6'h00;
      write_address_data_log_force[6591] <= 6'h00;
      write_address_data_log_force[6592] <= 6'h00;
      write_address_data_log_force[6593] <= 6'h00;
      write_address_data_log_force[6594] <= 6'h00;
      write_address_data_log_force[6595] <= 6'h00;
      write_address_data_log_force[6596] <= 6'h00;
      write_address_data_log_force[6597] <= 6'h00;
      write_address_data_log_force[6598] <= 6'h00;
      write_address_data_log_force[6599] <= 6'h00;
      write_address_data_log_force[6600] <= 6'h00;
      write_address_data_log_force[6601] <= 6'h00;
      write_address_data_log_force[6602] <= 6'h00;
      write_address_data_log_force[6603] <= 6'h00;
      write_address_data_log_force[6604] <= 6'h00;
      write_address_data_log_force[6605] <= 6'h00;
      write_address_data_log_force[6606] <= 6'h00;
      write_address_data_log_force[6607] <= 6'h00;
      write_address_data_log_force[6608] <= 6'h00;
      write_address_data_log_force[6609] <= 6'h00;
      write_address_data_log_force[6610] <= 6'h00;
      write_address_data_log_force[6611] <= 6'h00;
      write_address_data_log_force[6612] <= 6'h00;
      write_address_data_log_force[6613] <= 6'h00;
      write_address_data_log_force[6614] <= 6'h00;
      write_address_data_log_force[6615] <= 6'h00;
      write_address_data_log_force[6616] <= 6'h00;
      write_address_data_log_force[6617] <= 6'h00;
      write_address_data_log_force[6618] <= 6'h00;
      write_address_data_log_force[6619] <= 6'h00;
      write_address_data_log_force[6620] <= 6'h00;
      write_address_data_log_force[6621] <= 6'h00;
      write_address_data_log_force[6622] <= 6'h00;
      write_address_data_log_force[6623] <= 6'h00;
      write_address_data_log_force[6624] <= 6'h00;
      write_address_data_log_force[6625] <= 6'h00;
      write_address_data_log_force[6626] <= 6'h00;
      write_address_data_log_force[6627] <= 6'h00;
      write_address_data_log_force[6628] <= 6'h00;
      write_address_data_log_force[6629] <= 6'h00;
      write_address_data_log_force[6630] <= 6'h00;
      write_address_data_log_force[6631] <= 6'h00;
      write_address_data_log_force[6632] <= 6'h00;
      write_address_data_log_force[6633] <= 6'h00;
      write_address_data_log_force[6634] <= 6'h00;
      write_address_data_log_force[6635] <= 6'h00;
      write_address_data_log_force[6636] <= 6'h00;
      write_address_data_log_force[6637] <= 6'h00;
      write_address_data_log_force[6638] <= 6'h00;
      write_address_data_log_force[6639] <= 6'h00;
      write_address_data_log_force[6640] <= 6'h00;
      write_address_data_log_force[6641] <= 6'h00;
      write_address_data_log_force[6642] <= 6'h00;
      write_address_data_log_force[6643] <= 6'h00;
      write_address_data_log_force[6644] <= 6'h00;
      write_address_data_log_force[6645] <= 6'h00;
      write_address_data_log_force[6646] <= 6'h00;
      write_address_data_log_force[6647] <= 6'h00;
      write_address_data_log_force[6648] <= 6'h00;
      write_address_data_log_force[6649] <= 6'h00;
      write_address_data_log_force[6650] <= 6'h00;
      write_address_data_log_force[6651] <= 6'h00;
      write_address_data_log_force[6652] <= 6'h00;
      write_address_data_log_force[6653] <= 6'h00;
      write_address_data_log_force[6654] <= 6'h00;
      write_address_data_log_force[6655] <= 6'h00;
      write_address_data_log_force[6656] <= 6'h00;
      write_address_data_log_force[6657] <= 6'h00;
      write_address_data_log_force[6658] <= 6'h00;
      write_address_data_log_force[6659] <= 6'h00;
      write_address_data_log_force[6660] <= 6'h00;
      write_address_data_log_force[6661] <= 6'h00;
      write_address_data_log_force[6662] <= 6'h00;
      write_address_data_log_force[6663] <= 6'h00;
      write_address_data_log_force[6664] <= 6'h00;
      write_address_data_log_force[6665] <= 6'h00;
      write_address_data_log_force[6666] <= 6'h00;
      write_address_data_log_force[6667] <= 6'h00;
      write_address_data_log_force[6668] <= 6'h00;
      write_address_data_log_force[6669] <= 6'h00;
      write_address_data_log_force[6670] <= 6'h00;
      write_address_data_log_force[6671] <= 6'h00;
      write_address_data_log_force[6672] <= 6'h00;
      write_address_data_log_force[6673] <= 6'h00;
      write_address_data_log_force[6674] <= 6'h00;
      write_address_data_log_force[6675] <= 6'h00;
      write_address_data_log_force[6676] <= 6'h00;
      write_address_data_log_force[6677] <= 6'h00;
      write_address_data_log_force[6678] <= 6'h00;
      write_address_data_log_force[6679] <= 6'h00;
      write_address_data_log_force[6680] <= 6'h00;
      write_address_data_log_force[6681] <= 6'h00;
      write_address_data_log_force[6682] <= 6'h00;
      write_address_data_log_force[6683] <= 6'h00;
      write_address_data_log_force[6684] <= 6'h00;
      write_address_data_log_force[6685] <= 6'h00;
      write_address_data_log_force[6686] <= 6'h00;
      write_address_data_log_force[6687] <= 6'h00;
      write_address_data_log_force[6688] <= 6'h00;
      write_address_data_log_force[6689] <= 6'h00;
      write_address_data_log_force[6690] <= 6'h00;
      write_address_data_log_force[6691] <= 6'h00;
      write_address_data_log_force[6692] <= 6'h00;
      write_address_data_log_force[6693] <= 6'h00;
      write_address_data_log_force[6694] <= 6'h00;
      write_address_data_log_force[6695] <= 6'h00;
      write_address_data_log_force[6696] <= 6'h00;
      write_address_data_log_force[6697] <= 6'h00;
      write_address_data_log_force[6698] <= 6'h00;
      write_address_data_log_force[6699] <= 6'h00;
      write_address_data_log_force[6700] <= 6'h00;
      write_address_data_log_force[6701] <= 6'h00;
      write_address_data_log_force[6702] <= 6'h00;
      write_address_data_log_force[6703] <= 6'h00;
      write_address_data_log_force[6704] <= 6'h00;
      write_address_data_log_force[6705] <= 6'h00;
      write_address_data_log_force[6706] <= 6'h00;
      write_address_data_log_force[6707] <= 6'h00;
      write_address_data_log_force[6708] <= 6'h00;
      write_address_data_log_force[6709] <= 6'h00;
      write_address_data_log_force[6710] <= 6'h00;
      write_address_data_log_force[6711] <= 6'h00;
      write_address_data_log_force[6712] <= 6'h00;
      write_address_data_log_force[6713] <= 6'h00;
      write_address_data_log_force[6714] <= 6'h00;
      write_address_data_log_force[6715] <= 6'h00;
      write_address_data_log_force[6716] <= 6'h00;
      write_address_data_log_force[6717] <= 6'h00;
      write_address_data_log_force[6718] <= 6'h00;
      write_address_data_log_force[6719] <= 6'h00;
      write_address_data_log_force[6720] <= 6'h00;
      write_address_data_log_force[6721] <= 6'h00;
      write_address_data_log_force[6722] <= 6'h00;
      write_address_data_log_force[6723] <= 6'h00;
      write_address_data_log_force[6724] <= 6'h00;
      write_address_data_log_force[6725] <= 6'h00;
      write_address_data_log_force[6726] <= 6'h00;
      write_address_data_log_force[6727] <= 6'h00;
      write_address_data_log_force[6728] <= 6'h00;
      write_address_data_log_force[6729] <= 6'h00;
      write_address_data_log_force[6730] <= 6'h00;
      write_address_data_log_force[6731] <= 6'h00;
      write_address_data_log_force[6732] <= 6'h00;
      write_address_data_log_force[6733] <= 6'h00;
      write_address_data_log_force[6734] <= 6'h00;
      write_address_data_log_force[6735] <= 6'h00;
      write_address_data_log_force[6736] <= 6'h00;
      write_address_data_log_force[6737] <= 6'h00;
      write_address_data_log_force[6738] <= 6'h00;
      write_address_data_log_force[6739] <= 6'h00;
      write_address_data_log_force[6740] <= 6'h00;
      write_address_data_log_force[6741] <= 6'h00;
      write_address_data_log_force[6742] <= 6'h00;
      write_address_data_log_force[6743] <= 6'h00;
      write_address_data_log_force[6744] <= 6'h00;
      write_address_data_log_force[6745] <= 6'h00;
      write_address_data_log_force[6746] <= 6'h00;
      write_address_data_log_force[6747] <= 6'h00;
      write_address_data_log_force[6748] <= 6'h00;
      write_address_data_log_force[6749] <= 6'h00;
      write_address_data_log_force[6750] <= 6'h00;
      write_address_data_log_force[6751] <= 6'h00;
      write_address_data_log_force[6752] <= 6'h00;
      write_address_data_log_force[6753] <= 6'h00;
      write_address_data_log_force[6754] <= 6'h00;
      write_address_data_log_force[6755] <= 6'h00;
      write_address_data_log_force[6756] <= 6'h00;
      write_address_data_log_force[6757] <= 6'h00;
      write_address_data_log_force[6758] <= 6'h00;
      write_address_data_log_force[6759] <= 6'h00;
      write_address_data_log_force[6760] <= 6'h00;
      write_address_data_log_force[6761] <= 6'h00;
      write_address_data_log_force[6762] <= 6'h00;
      write_address_data_log_force[6763] <= 6'h00;
      write_address_data_log_force[6764] <= 6'h00;
      write_address_data_log_force[6765] <= 6'h00;
      write_address_data_log_force[6766] <= 6'h00;
      write_address_data_log_force[6767] <= 6'h00;
      write_address_data_log_force[6768] <= 6'h00;
      write_address_data_log_force[6769] <= 6'h00;
      write_address_data_log_force[6770] <= 6'h00;
      write_address_data_log_force[6771] <= 6'h00;
      write_address_data_log_force[6772] <= 6'h00;
      write_address_data_log_force[6773] <= 6'h00;
      write_address_data_log_force[6774] <= 6'h00;
      write_address_data_log_force[6775] <= 6'h00;
      write_address_data_log_force[6776] <= 6'h00;
      write_address_data_log_force[6777] <= 6'h00;
      write_address_data_log_force[6778] <= 6'h00;
      write_address_data_log_force[6779] <= 6'h00;
      write_address_data_log_force[6780] <= 6'h00;
      write_address_data_log_force[6781] <= 6'h00;
      write_address_data_log_force[6782] <= 6'h00;
      write_address_data_log_force[6783] <= 6'h00;
      write_address_data_log_force[6784] <= 6'h00;
      write_address_data_log_force[6785] <= 6'h00;
      write_address_data_log_force[6786] <= 6'h00;
      write_address_data_log_force[6787] <= 6'h00;
      write_address_data_log_force[6788] <= 6'h00;
      write_address_data_log_force[6789] <= 6'h00;
      write_address_data_log_force[6790] <= 6'h00;
      write_address_data_log_force[6791] <= 6'h00;
      write_address_data_log_force[6792] <= 6'h00;
      write_address_data_log_force[6793] <= 6'h00;
      write_address_data_log_force[6794] <= 6'h00;
      write_address_data_log_force[6795] <= 6'h00;
      write_address_data_log_force[6796] <= 6'h00;
      write_address_data_log_force[6797] <= 6'h00;
      write_address_data_log_force[6798] <= 6'h00;
      write_address_data_log_force[6799] <= 6'h00;
      write_address_data_log_force[6800] <= 6'h00;
      write_address_data_log_force[6801] <= 6'h00;
      write_address_data_log_force[6802] <= 6'h00;
      write_address_data_log_force[6803] <= 6'h00;
      write_address_data_log_force[6804] <= 6'h00;
      write_address_data_log_force[6805] <= 6'h00;
      write_address_data_log_force[6806] <= 6'h00;
      write_address_data_log_force[6807] <= 6'h00;
      write_address_data_log_force[6808] <= 6'h00;
      write_address_data_log_force[6809] <= 6'h00;
      write_address_data_log_force[6810] <= 6'h00;
      write_address_data_log_force[6811] <= 6'h00;
      write_address_data_log_force[6812] <= 6'h00;
      write_address_data_log_force[6813] <= 6'h00;
      write_address_data_log_force[6814] <= 6'h00;
      write_address_data_log_force[6815] <= 6'h00;
      write_address_data_log_force[6816] <= 6'h00;
      write_address_data_log_force[6817] <= 6'h00;
      write_address_data_log_force[6818] <= 6'h00;
      write_address_data_log_force[6819] <= 6'h00;
      write_address_data_log_force[6820] <= 6'h00;
      write_address_data_log_force[6821] <= 6'h00;
      write_address_data_log_force[6822] <= 6'h00;
      write_address_data_log_force[6823] <= 6'h00;
      write_address_data_log_force[6824] <= 6'h00;
      write_address_data_log_force[6825] <= 6'h00;
      write_address_data_log_force[6826] <= 6'h00;
      write_address_data_log_force[6827] <= 6'h00;
      write_address_data_log_force[6828] <= 6'h00;
      write_address_data_log_force[6829] <= 6'h00;
      write_address_data_log_force[6830] <= 6'h00;
      write_address_data_log_force[6831] <= 6'h00;
      write_address_data_log_force[6832] <= 6'h00;
      write_address_data_log_force[6833] <= 6'h00;
      write_address_data_log_force[6834] <= 6'h00;
      write_address_data_log_force[6835] <= 6'h00;
      write_address_data_log_force[6836] <= 6'h00;
      write_address_data_log_force[6837] <= 6'h00;
      write_address_data_log_force[6838] <= 6'h00;
      write_address_data_log_force[6839] <= 6'h00;
      write_address_data_log_force[6840] <= 6'h00;
      write_address_data_log_force[6841] <= 6'h00;
      write_address_data_log_force[6842] <= 6'h00;
      write_address_data_log_force[6843] <= 6'h00;
      write_address_data_log_force[6844] <= 6'h00;
      write_address_data_log_force[6845] <= 6'h00;
      write_address_data_log_force[6846] <= 6'h00;
      write_address_data_log_force[6847] <= 6'h00;
      write_address_data_log_force[6848] <= 6'h00;
      write_address_data_log_force[6849] <= 6'h00;
      write_address_data_log_force[6850] <= 6'h00;
      write_address_data_log_force[6851] <= 6'h00;
      write_address_data_log_force[6852] <= 6'h00;
      write_address_data_log_force[6853] <= 6'h00;
      write_address_data_log_force[6854] <= 6'h00;
      write_address_data_log_force[6855] <= 6'h00;
      write_address_data_log_force[6856] <= 6'h00;
      write_address_data_log_force[6857] <= 6'h00;
      write_address_data_log_force[6858] <= 6'h00;
      write_address_data_log_force[6859] <= 6'h00;
      write_address_data_log_force[6860] <= 6'h00;
      write_address_data_log_force[6861] <= 6'h00;
      write_address_data_log_force[6862] <= 6'h00;
      write_address_data_log_force[6863] <= 6'h00;
      write_address_data_log_force[6864] <= 6'h00;
      write_address_data_log_force[6865] <= 6'h00;
      write_address_data_log_force[6866] <= 6'h00;
      write_address_data_log_force[6867] <= 6'h00;
      write_address_data_log_force[6868] <= 6'h00;
      write_address_data_log_force[6869] <= 6'h00;
      write_address_data_log_force[6870] <= 6'h00;
      write_address_data_log_force[6871] <= 6'h00;
      write_address_data_log_force[6872] <= 6'h00;
      write_address_data_log_force[6873] <= 6'h00;
      write_address_data_log_force[6874] <= 6'h00;
      write_address_data_log_force[6875] <= 6'h00;
      write_address_data_log_force[6876] <= 6'h00;
      write_address_data_log_force[6877] <= 6'h00;
      write_address_data_log_force[6878] <= 6'h00;
      write_address_data_log_force[6879] <= 6'h00;
      write_address_data_log_force[6880] <= 6'h00;
      write_address_data_log_force[6881] <= 6'h00;
      write_address_data_log_force[6882] <= 6'h00;
      write_address_data_log_force[6883] <= 6'h00;
      write_address_data_log_force[6884] <= 6'h00;
      write_address_data_log_force[6885] <= 6'h00;
      write_address_data_log_force[6886] <= 6'h00;
      write_address_data_log_force[6887] <= 6'h00;
      write_address_data_log_force[6888] <= 6'h00;
      write_address_data_log_force[6889] <= 6'h00;
      write_address_data_log_force[6890] <= 6'h00;
      write_address_data_log_force[6891] <= 6'h00;
      write_address_data_log_force[6892] <= 6'h00;
      write_address_data_log_force[6893] <= 6'h00;
      write_address_data_log_force[6894] <= 6'h00;
      write_address_data_log_force[6895] <= 6'h00;
      write_address_data_log_force[6896] <= 6'h00;
      write_address_data_log_force[6897] <= 6'h00;
      write_address_data_log_force[6898] <= 6'h00;
      write_address_data_log_force[6899] <= 6'h00;
      write_address_data_log_force[6900] <= 6'h00;
      write_address_data_log_force[6901] <= 6'h00;
      write_address_data_log_force[6902] <= 6'h00;
      write_address_data_log_force[6903] <= 6'h00;
      write_address_data_log_force[6904] <= 6'h00;
      write_address_data_log_force[6905] <= 6'h00;
      write_address_data_log_force[6906] <= 6'h00;
      write_address_data_log_force[6907] <= 6'h00;
      write_address_data_log_force[6908] <= 6'h00;
      write_address_data_log_force[6909] <= 6'h00;
      write_address_data_log_force[6910] <= 6'h00;
      write_address_data_log_force[6911] <= 6'h00;
      write_address_data_log_force[6912] <= 6'h00;
      write_address_data_log_force[6913] <= 6'h00;
      write_address_data_log_force[6914] <= 6'h00;
      write_address_data_log_force[6915] <= 6'h00;
      write_address_data_log_force[6916] <= 6'h00;
      write_address_data_log_force[6917] <= 6'h00;
      write_address_data_log_force[6918] <= 6'h00;
      write_address_data_log_force[6919] <= 6'h00;
      write_address_data_log_force[6920] <= 6'h00;
      write_address_data_log_force[6921] <= 6'h00;
      write_address_data_log_force[6922] <= 6'h00;
      write_address_data_log_force[6923] <= 6'h00;
      write_address_data_log_force[6924] <= 6'h00;
      write_address_data_log_force[6925] <= 6'h00;
      write_address_data_log_force[6926] <= 6'h00;
      write_address_data_log_force[6927] <= 6'h00;
      write_address_data_log_force[6928] <= 6'h00;
      write_address_data_log_force[6929] <= 6'h00;
      write_address_data_log_force[6930] <= 6'h00;
      write_address_data_log_force[6931] <= 6'h00;
      write_address_data_log_force[6932] <= 6'h00;
      write_address_data_log_force[6933] <= 6'h00;
      write_address_data_log_force[6934] <= 6'h00;
      write_address_data_log_force[6935] <= 6'h00;
      write_address_data_log_force[6936] <= 6'h00;
      write_address_data_log_force[6937] <= 6'h00;
      write_address_data_log_force[6938] <= 6'h00;
      write_address_data_log_force[6939] <= 6'h00;
      write_address_data_log_force[6940] <= 6'h00;
      write_address_data_log_force[6941] <= 6'h00;
      write_address_data_log_force[6942] <= 6'h00;
      write_address_data_log_force[6943] <= 6'h00;
      write_address_data_log_force[6944] <= 6'h00;
      write_address_data_log_force[6945] <= 6'h00;
      write_address_data_log_force[6946] <= 6'h00;
      write_address_data_log_force[6947] <= 6'h00;
      write_address_data_log_force[6948] <= 6'h00;
      write_address_data_log_force[6949] <= 6'h00;
      write_address_data_log_force[6950] <= 6'h00;
      write_address_data_log_force[6951] <= 6'h00;
      write_address_data_log_force[6952] <= 6'h00;
      write_address_data_log_force[6953] <= 6'h00;
      write_address_data_log_force[6954] <= 6'h00;
      write_address_data_log_force[6955] <= 6'h00;
      write_address_data_log_force[6956] <= 6'h00;
      write_address_data_log_force[6957] <= 6'h00;
      write_address_data_log_force[6958] <= 6'h00;
      write_address_data_log_force[6959] <= 6'h00;
      write_address_data_log_force[6960] <= 6'h00;
      write_address_data_log_force[6961] <= 6'h00;
      write_address_data_log_force[6962] <= 6'h00;
      write_address_data_log_force[6963] <= 6'h00;
      write_address_data_log_force[6964] <= 6'h00;
      write_address_data_log_force[6965] <= 6'h00;
      write_address_data_log_force[6966] <= 6'h00;
      write_address_data_log_force[6967] <= 6'h00;
      write_address_data_log_force[6968] <= 6'h00;
      write_address_data_log_force[6969] <= 6'h00;
      write_address_data_log_force[6970] <= 6'h00;
      write_address_data_log_force[6971] <= 6'h00;
      write_address_data_log_force[6972] <= 6'h00;
      write_address_data_log_force[6973] <= 6'h00;
      write_address_data_log_force[6974] <= 6'h00;
      write_address_data_log_force[6975] <= 6'h00;
      write_address_data_log_force[6976] <= 6'h00;
      write_address_data_log_force[6977] <= 6'h00;
      write_address_data_log_force[6978] <= 6'h00;
      write_address_data_log_force[6979] <= 6'h00;
      write_address_data_log_force[6980] <= 6'h00;
      write_address_data_log_force[6981] <= 6'h00;
      write_address_data_log_force[6982] <= 6'h00;
      write_address_data_log_force[6983] <= 6'h00;
      write_address_data_log_force[6984] <= 6'h00;
      write_address_data_log_force[6985] <= 6'h00;
      write_address_data_log_force[6986] <= 6'h00;
      write_address_data_log_force[6987] <= 6'h00;
      write_address_data_log_force[6988] <= 6'h00;
      write_address_data_log_force[6989] <= 6'h00;
      write_address_data_log_force[6990] <= 6'h00;
      write_address_data_log_force[6991] <= 6'h00;
      write_address_data_log_force[6992] <= 6'h00;
      write_address_data_log_force[6993] <= 6'h00;
      write_address_data_log_force[6994] <= 6'h00;
      write_address_data_log_force[6995] <= 6'h00;
      write_address_data_log_force[6996] <= 6'h00;
      write_address_data_log_force[6997] <= 6'h00;
      write_address_data_log_force[6998] <= 6'h00;
      write_address_data_log_force[6999] <= 6'h00;
      write_address_data_log_force[7000] <= 6'h00;
      write_address_data_log_force[7001] <= 6'h00;
      write_address_data_log_force[7002] <= 6'h00;
      write_address_data_log_force[7003] <= 6'h00;
      write_address_data_log_force[7004] <= 6'h00;
      write_address_data_log_force[7005] <= 6'h00;
      write_address_data_log_force[7006] <= 6'h00;
      write_address_data_log_force[7007] <= 6'h00;
      write_address_data_log_force[7008] <= 6'h00;
      write_address_data_log_force[7009] <= 6'h00;
      write_address_data_log_force[7010] <= 6'h00;
      write_address_data_log_force[7011] <= 6'h00;
      write_address_data_log_force[7012] <= 6'h00;
      write_address_data_log_force[7013] <= 6'h00;
      write_address_data_log_force[7014] <= 6'h00;
      write_address_data_log_force[7015] <= 6'h00;
      write_address_data_log_force[7016] <= 6'h00;
      write_address_data_log_force[7017] <= 6'h00;
      write_address_data_log_force[7018] <= 6'h00;
      write_address_data_log_force[7019] <= 6'h00;
      write_address_data_log_force[7020] <= 6'h00;
      write_address_data_log_force[7021] <= 6'h00;
      write_address_data_log_force[7022] <= 6'h00;
      write_address_data_log_force[7023] <= 6'h00;
      write_address_data_log_force[7024] <= 6'h00;
      write_address_data_log_force[7025] <= 6'h00;
      write_address_data_log_force[7026] <= 6'h00;
      write_address_data_log_force[7027] <= 6'h00;
      write_address_data_log_force[7028] <= 6'h00;
      write_address_data_log_force[7029] <= 6'h00;
      write_address_data_log_force[7030] <= 6'h00;
      write_address_data_log_force[7031] <= 6'h00;
      write_address_data_log_force[7032] <= 6'h00;
      write_address_data_log_force[7033] <= 6'h00;
      write_address_data_log_force[7034] <= 6'h00;
      write_address_data_log_force[7035] <= 6'h00;
      write_address_data_log_force[7036] <= 6'h00;
      write_address_data_log_force[7037] <= 6'h00;
      write_address_data_log_force[7038] <= 6'h00;
      write_address_data_log_force[7039] <= 6'h00;
      write_address_data_log_force[7040] <= 6'h00;
      write_address_data_log_force[7041] <= 6'h00;
      write_address_data_log_force[7042] <= 6'h00;
      write_address_data_log_force[7043] <= 6'h00;
      write_address_data_log_force[7044] <= 6'h00;
      write_address_data_log_force[7045] <= 6'h00;
      write_address_data_log_force[7046] <= 6'h00;
      write_address_data_log_force[7047] <= 6'h00;
      write_address_data_log_force[7048] <= 6'h00;
      write_address_data_log_force[7049] <= 6'h00;
      write_address_data_log_force[7050] <= 6'h00;
      write_address_data_log_force[7051] <= 6'h00;
      write_address_data_log_force[7052] <= 6'h00;
      write_address_data_log_force[7053] <= 6'h00;
      write_address_data_log_force[7054] <= 6'h00;
      write_address_data_log_force[7055] <= 6'h00;
      write_address_data_log_force[7056] <= 6'h00;
      write_address_data_log_force[7057] <= 6'h00;
      write_address_data_log_force[7058] <= 6'h00;
      write_address_data_log_force[7059] <= 6'h00;
      write_address_data_log_force[7060] <= 6'h00;
      write_address_data_log_force[7061] <= 6'h00;
      write_address_data_log_force[7062] <= 6'h00;
      write_address_data_log_force[7063] <= 6'h00;
      write_address_data_log_force[7064] <= 6'h00;
      write_address_data_log_force[7065] <= 6'h00;
      write_address_data_log_force[7066] <= 6'h00;
      write_address_data_log_force[7067] <= 6'h00;
      write_address_data_log_force[7068] <= 6'h00;
      write_address_data_log_force[7069] <= 6'h00;
      write_address_data_log_force[7070] <= 6'h00;
      write_address_data_log_force[7071] <= 6'h00;
      write_address_data_log_force[7072] <= 6'h00;
      write_address_data_log_force[7073] <= 6'h00;
      write_address_data_log_force[7074] <= 6'h00;
      write_address_data_log_force[7075] <= 6'h00;
      write_address_data_log_force[7076] <= 6'h00;
      write_address_data_log_force[7077] <= 6'h00;
      write_address_data_log_force[7078] <= 6'h00;
      write_address_data_log_force[7079] <= 6'h00;
      write_address_data_log_force[7080] <= 6'h00;
      write_address_data_log_force[7081] <= 6'h00;
      write_address_data_log_force[7082] <= 6'h00;
      write_address_data_log_force[7083] <= 6'h00;
      write_address_data_log_force[7084] <= 6'h00;
      write_address_data_log_force[7085] <= 6'h00;
      write_address_data_log_force[7086] <= 6'h00;
      write_address_data_log_force[7087] <= 6'h00;
      write_address_data_log_force[7088] <= 6'h00;
      write_address_data_log_force[7089] <= 6'h00;
      write_address_data_log_force[7090] <= 6'h00;
      write_address_data_log_force[7091] <= 6'h00;
      write_address_data_log_force[7092] <= 6'h00;
      write_address_data_log_force[7093] <= 6'h00;
      write_address_data_log_force[7094] <= 6'h00;
      write_address_data_log_force[7095] <= 6'h00;
      write_address_data_log_force[7096] <= 6'h00;
      write_address_data_log_force[7097] <= 6'h00;
      write_address_data_log_force[7098] <= 6'h00;
      write_address_data_log_force[7099] <= 6'h00;
      write_address_data_log_force[7100] <= 6'h00;
      write_address_data_log_force[7101] <= 6'h00;
      write_address_data_log_force[7102] <= 6'h00;
      write_address_data_log_force[7103] <= 6'h00;
      write_address_data_log_force[7104] <= 6'h00;
      write_address_data_log_force[7105] <= 6'h00;
      write_address_data_log_force[7106] <= 6'h00;
      write_address_data_log_force[7107] <= 6'h00;
      write_address_data_log_force[7108] <= 6'h00;
      write_address_data_log_force[7109] <= 6'h00;
      write_address_data_log_force[7110] <= 6'h00;
      write_address_data_log_force[7111] <= 6'h00;
      write_address_data_log_force[7112] <= 6'h00;
      write_address_data_log_force[7113] <= 6'h00;
      write_address_data_log_force[7114] <= 6'h00;
      write_address_data_log_force[7115] <= 6'h00;
      write_address_data_log_force[7116] <= 6'h00;
      write_address_data_log_force[7117] <= 6'h00;
      write_address_data_log_force[7118] <= 6'h00;
      write_address_data_log_force[7119] <= 6'h00;
      write_address_data_log_force[7120] <= 6'h00;
      write_address_data_log_force[7121] <= 6'h00;
      write_address_data_log_force[7122] <= 6'h00;
      write_address_data_log_force[7123] <= 6'h00;
      write_address_data_log_force[7124] <= 6'h00;
      write_address_data_log_force[7125] <= 6'h00;
      write_address_data_log_force[7126] <= 6'h00;
      write_address_data_log_force[7127] <= 6'h00;
      write_address_data_log_force[7128] <= 6'h00;
      write_address_data_log_force[7129] <= 6'h00;
      write_address_data_log_force[7130] <= 6'h00;
      write_address_data_log_force[7131] <= 6'h00;
      write_address_data_log_force[7132] <= 6'h00;
      write_address_data_log_force[7133] <= 6'h00;
      write_address_data_log_force[7134] <= 6'h00;
      write_address_data_log_force[7135] <= 6'h00;
      write_address_data_log_force[7136] <= 6'h00;
      write_address_data_log_force[7137] <= 6'h00;
      write_address_data_log_force[7138] <= 6'h00;
      write_address_data_log_force[7139] <= 6'h00;
      write_address_data_log_force[7140] <= 6'h00;
      write_address_data_log_force[7141] <= 6'h00;
      write_address_data_log_force[7142] <= 6'h00;
      write_address_data_log_force[7143] <= 6'h00;
      write_address_data_log_force[7144] <= 6'h00;
      write_address_data_log_force[7145] <= 6'h00;
      write_address_data_log_force[7146] <= 6'h00;
      write_address_data_log_force[7147] <= 6'h00;
      write_address_data_log_force[7148] <= 6'h00;
      write_address_data_log_force[7149] <= 6'h00;
      write_address_data_log_force[7150] <= 6'h00;
      write_address_data_log_force[7151] <= 6'h00;
      write_address_data_log_force[7152] <= 6'h00;
      write_address_data_log_force[7153] <= 6'h00;
      write_address_data_log_force[7154] <= 6'h00;
      write_address_data_log_force[7155] <= 6'h00;
      write_address_data_log_force[7156] <= 6'h00;
      write_address_data_log_force[7157] <= 6'h00;
      write_address_data_log_force[7158] <= 6'h00;
      write_address_data_log_force[7159] <= 6'h00;
      write_address_data_log_force[7160] <= 6'h00;
      write_address_data_log_force[7161] <= 6'h00;
      write_address_data_log_force[7162] <= 6'h00;
      write_address_data_log_force[7163] <= 6'h00;
      write_address_data_log_force[7164] <= 6'h00;
      write_address_data_log_force[7165] <= 6'h00;
      write_address_data_log_force[7166] <= 6'h00;
      write_address_data_log_force[7167] <= 6'h00;
      write_address_data_log_force[7168] <= 6'h00;
      write_address_data_log_force[7169] <= 6'h00;
      write_address_data_log_force[7170] <= 6'h00;
      write_address_data_log_force[7171] <= 6'h00;
      write_address_data_log_force[7172] <= 6'h00;
      write_address_data_log_force[7173] <= 6'h00;
      write_address_data_log_force[7174] <= 6'h00;
      write_address_data_log_force[7175] <= 6'h00;
      write_address_data_log_force[7176] <= 6'h00;
      write_address_data_log_force[7177] <= 6'h00;
      write_address_data_log_force[7178] <= 6'h00;
      write_address_data_log_force[7179] <= 6'h00;
      write_address_data_log_force[7180] <= 6'h00;
      write_address_data_log_force[7181] <= 6'h00;
      write_address_data_log_force[7182] <= 6'h00;
      write_address_data_log_force[7183] <= 6'h00;
      write_address_data_log_force[7184] <= 6'h00;
      write_address_data_log_force[7185] <= 6'h00;
      write_address_data_log_force[7186] <= 6'h00;
      write_address_data_log_force[7187] <= 6'h00;
      write_address_data_log_force[7188] <= 6'h00;
      write_address_data_log_force[7189] <= 6'h00;
      write_address_data_log_force[7190] <= 6'h00;
      write_address_data_log_force[7191] <= 6'h00;
      write_address_data_log_force[7192] <= 6'h00;
      write_address_data_log_force[7193] <= 6'h00;
      write_address_data_log_force[7194] <= 6'h00;
      write_address_data_log_force[7195] <= 6'h00;
      write_address_data_log_force[7196] <= 6'h00;
      write_address_data_log_force[7197] <= 6'h00;
      write_address_data_log_force[7198] <= 6'h00;
      write_address_data_log_force[7199] <= 6'h00;
      write_address_data_log_force[7200] <= 6'h00;
      write_address_data_log_force[7201] <= 6'h00;
      write_address_data_log_force[7202] <= 6'h00;
      write_address_data_log_force[7203] <= 6'h00;
      write_address_data_log_force[7204] <= 6'h00;
      write_address_data_log_force[7205] <= 6'h00;
      write_address_data_log_force[7206] <= 6'h00;
      write_address_data_log_force[7207] <= 6'h00;
      write_address_data_log_force[7208] <= 6'h00;
      write_address_data_log_force[7209] <= 6'h00;
      write_address_data_log_force[7210] <= 6'h00;
      write_address_data_log_force[7211] <= 6'h00;
      write_address_data_log_force[7212] <= 6'h00;
      write_address_data_log_force[7213] <= 6'h00;
      write_address_data_log_force[7214] <= 6'h00;
      write_address_data_log_force[7215] <= 6'h00;
      write_address_data_log_force[7216] <= 6'h00;
      write_address_data_log_force[7217] <= 6'h00;
      write_address_data_log_force[7218] <= 6'h00;
      write_address_data_log_force[7219] <= 6'h00;
      write_address_data_log_force[7220] <= 6'h00;
      write_address_data_log_force[7221] <= 6'h00;
      write_address_data_log_force[7222] <= 6'h00;
      write_address_data_log_force[7223] <= 6'h00;
      write_address_data_log_force[7224] <= 6'h00;
      write_address_data_log_force[7225] <= 6'h00;
      write_address_data_log_force[7226] <= 6'h00;
      write_address_data_log_force[7227] <= 6'h00;
      write_address_data_log_force[7228] <= 6'h00;
      write_address_data_log_force[7229] <= 6'h00;
      write_address_data_log_force[7230] <= 6'h00;
      write_address_data_log_force[7231] <= 6'h00;
      write_address_data_log_force[7232] <= 6'h00;
      write_address_data_log_force[7233] <= 6'h00;
      write_address_data_log_force[7234] <= 6'h00;
      write_address_data_log_force[7235] <= 6'h00;
      write_address_data_log_force[7236] <= 6'h00;
      write_address_data_log_force[7237] <= 6'h00;
      write_address_data_log_force[7238] <= 6'h00;
      write_address_data_log_force[7239] <= 6'h00;
      write_address_data_log_force[7240] <= 6'h00;
      write_address_data_log_force[7241] <= 6'h00;
      write_address_data_log_force[7242] <= 6'h00;
      write_address_data_log_force[7243] <= 6'h00;
      write_address_data_log_force[7244] <= 6'h00;
      write_address_data_log_force[7245] <= 6'h00;
      write_address_data_log_force[7246] <= 6'h00;
      write_address_data_log_force[7247] <= 6'h00;
      write_address_data_log_force[7248] <= 6'h00;
      write_address_data_log_force[7249] <= 6'h00;
      write_address_data_log_force[7250] <= 6'h00;
      write_address_data_log_force[7251] <= 6'h00;
      write_address_data_log_force[7252] <= 6'h00;
      write_address_data_log_force[7253] <= 6'h00;
      write_address_data_log_force[7254] <= 6'h00;
      write_address_data_log_force[7255] <= 6'h00;
      write_address_data_log_force[7256] <= 6'h00;
      write_address_data_log_force[7257] <= 6'h00;
      write_address_data_log_force[7258] <= 6'h00;
      write_address_data_log_force[7259] <= 6'h00;
      write_address_data_log_force[7260] <= 6'h00;
      write_address_data_log_force[7261] <= 6'h00;
      write_address_data_log_force[7262] <= 6'h00;
      write_address_data_log_force[7263] <= 6'h00;
      write_address_data_log_force[7264] <= 6'h00;
      write_address_data_log_force[7265] <= 6'h00;
      write_address_data_log_force[7266] <= 6'h00;
      write_address_data_log_force[7267] <= 6'h00;
      write_address_data_log_force[7268] <= 6'h00;
      write_address_data_log_force[7269] <= 6'h00;
      write_address_data_log_force[7270] <= 6'h00;
      write_address_data_log_force[7271] <= 6'h00;
      write_address_data_log_force[7272] <= 6'h00;
      write_address_data_log_force[7273] <= 6'h00;
      write_address_data_log_force[7274] <= 6'h00;
      write_address_data_log_force[7275] <= 6'h00;
      write_address_data_log_force[7276] <= 6'h00;
      write_address_data_log_force[7277] <= 6'h00;
      write_address_data_log_force[7278] <= 6'h00;
      write_address_data_log_force[7279] <= 6'h00;
      write_address_data_log_force[7280] <= 6'h00;
      write_address_data_log_force[7281] <= 6'h00;
      write_address_data_log_force[7282] <= 6'h00;
      write_address_data_log_force[7283] <= 6'h00;
      write_address_data_log_force[7284] <= 6'h00;
      write_address_data_log_force[7285] <= 6'h00;
      write_address_data_log_force[7286] <= 6'h00;
      write_address_data_log_force[7287] <= 6'h00;
      write_address_data_log_force[7288] <= 6'h00;
      write_address_data_log_force[7289] <= 6'h00;
      write_address_data_log_force[7290] <= 6'h00;
      write_address_data_log_force[7291] <= 6'h00;
      write_address_data_log_force[7292] <= 6'h00;
      write_address_data_log_force[7293] <= 6'h00;
      write_address_data_log_force[7294] <= 6'h00;
      write_address_data_log_force[7295] <= 6'h00;
      write_address_data_log_force[7296] <= 6'h00;
      write_address_data_log_force[7297] <= 6'h00;
      write_address_data_log_force[7298] <= 6'h00;
      write_address_data_log_force[7299] <= 6'h00;
      write_address_data_log_force[7300] <= 6'h00;
      write_address_data_log_force[7301] <= 6'h00;
      write_address_data_log_force[7302] <= 6'h00;
      write_address_data_log_force[7303] <= 6'h00;
      write_address_data_log_force[7304] <= 6'h00;
      write_address_data_log_force[7305] <= 6'h00;
      write_address_data_log_force[7306] <= 6'h00;
      write_address_data_log_force[7307] <= 6'h00;
      write_address_data_log_force[7308] <= 6'h00;
      write_address_data_log_force[7309] <= 6'h00;
      write_address_data_log_force[7310] <= 6'h00;
      write_address_data_log_force[7311] <= 6'h00;
      write_address_data_log_force[7312] <= 6'h00;
      write_address_data_log_force[7313] <= 6'h00;
      write_address_data_log_force[7314] <= 6'h00;
      write_address_data_log_force[7315] <= 6'h00;
      write_address_data_log_force[7316] <= 6'h00;
      write_address_data_log_force[7317] <= 6'h00;
      write_address_data_log_force[7318] <= 6'h00;
      write_address_data_log_force[7319] <= 6'h00;
      write_address_data_log_force[7320] <= 6'h00;
      write_address_data_log_force[7321] <= 6'h00;
      write_address_data_log_force[7322] <= 6'h00;
      write_address_data_log_force[7323] <= 6'h00;
      write_address_data_log_force[7324] <= 6'h00;
      write_address_data_log_force[7325] <= 6'h00;
      write_address_data_log_force[7326] <= 6'h00;
      write_address_data_log_force[7327] <= 6'h00;
      write_address_data_log_force[7328] <= 6'h00;
      write_address_data_log_force[7329] <= 6'h00;
      write_address_data_log_force[7330] <= 6'h00;
      write_address_data_log_force[7331] <= 6'h00;
      write_address_data_log_force[7332] <= 6'h00;
      write_address_data_log_force[7333] <= 6'h00;
      write_address_data_log_force[7334] <= 6'h00;
      write_address_data_log_force[7335] <= 6'h00;
      write_address_data_log_force[7336] <= 6'h00;
      write_address_data_log_force[7337] <= 6'h00;
      write_address_data_log_force[7338] <= 6'h00;
      write_address_data_log_force[7339] <= 6'h00;
      write_address_data_log_force[7340] <= 6'h00;
      write_address_data_log_force[7341] <= 6'h00;
      write_address_data_log_force[7342] <= 6'h00;
      write_address_data_log_force[7343] <= 6'h00;
      write_address_data_log_force[7344] <= 6'h00;
      write_address_data_log_force[7345] <= 6'h00;
      write_address_data_log_force[7346] <= 6'h00;
      write_address_data_log_force[7347] <= 6'h00;
      write_address_data_log_force[7348] <= 6'h00;
      write_address_data_log_force[7349] <= 6'h00;
      write_address_data_log_force[7350] <= 6'h00;
      write_address_data_log_force[7351] <= 6'h00;
      write_address_data_log_force[7352] <= 6'h00;
      write_address_data_log_force[7353] <= 6'h00;
      write_address_data_log_force[7354] <= 6'h00;
      write_address_data_log_force[7355] <= 6'h00;
      write_address_data_log_force[7356] <= 6'h00;
      write_address_data_log_force[7357] <= 6'h00;
      write_address_data_log_force[7358] <= 6'h00;
      write_address_data_log_force[7359] <= 6'h00;
      write_address_data_log_force[7360] <= 6'h00;
      write_address_data_log_force[7361] <= 6'h00;
      write_address_data_log_force[7362] <= 6'h00;
      write_address_data_log_force[7363] <= 6'h00;
      write_address_data_log_force[7364] <= 6'h00;
      write_address_data_log_force[7365] <= 6'h00;
      write_address_data_log_force[7366] <= 6'h00;
      write_address_data_log_force[7367] <= 6'h00;
      write_address_data_log_force[7368] <= 6'h00;
      write_address_data_log_force[7369] <= 6'h00;
      write_address_data_log_force[7370] <= 6'h00;
      write_address_data_log_force[7371] <= 6'h00;
      write_address_data_log_force[7372] <= 6'h00;
      write_address_data_log_force[7373] <= 6'h00;
      write_address_data_log_force[7374] <= 6'h00;
      write_address_data_log_force[7375] <= 6'h00;
      write_address_data_log_force[7376] <= 6'h00;
      write_address_data_log_force[7377] <= 6'h00;
      write_address_data_log_force[7378] <= 6'h00;
      write_address_data_log_force[7379] <= 6'h00;
      write_address_data_log_force[7380] <= 6'h00;
      write_address_data_log_force[7381] <= 6'h00;
      write_address_data_log_force[7382] <= 6'h00;
      write_address_data_log_force[7383] <= 6'h00;
      write_address_data_log_force[7384] <= 6'h00;
      write_address_data_log_force[7385] <= 6'h00;
      write_address_data_log_force[7386] <= 6'h00;
      write_address_data_log_force[7387] <= 6'h00;
      write_address_data_log_force[7388] <= 6'h00;
      write_address_data_log_force[7389] <= 6'h00;
      write_address_data_log_force[7390] <= 6'h00;
      write_address_data_log_force[7391] <= 6'h00;
      write_address_data_log_force[7392] <= 6'h00;
      write_address_data_log_force[7393] <= 6'h00;
      write_address_data_log_force[7394] <= 6'h00;
      write_address_data_log_force[7395] <= 6'h00;
      write_address_data_log_force[7396] <= 6'h00;
      write_address_data_log_force[7397] <= 6'h00;
      write_address_data_log_force[7398] <= 6'h00;
      write_address_data_log_force[7399] <= 6'h00;
      write_address_data_log_force[7400] <= 6'h00;
      write_address_data_log_force[7401] <= 6'h00;
      write_address_data_log_force[7402] <= 6'h00;
      write_address_data_log_force[7403] <= 6'h00;
      write_address_data_log_force[7404] <= 6'h00;
      write_address_data_log_force[7405] <= 6'h00;
      write_address_data_log_force[7406] <= 6'h00;
      write_address_data_log_force[7407] <= 6'h00;
      write_address_data_log_force[7408] <= 6'h00;
      write_address_data_log_force[7409] <= 6'h00;
      write_address_data_log_force[7410] <= 6'h00;
      write_address_data_log_force[7411] <= 6'h00;
      write_address_data_log_force[7412] <= 6'h00;
      write_address_data_log_force[7413] <= 6'h00;
      write_address_data_log_force[7414] <= 6'h00;
      write_address_data_log_force[7415] <= 6'h00;
      write_address_data_log_force[7416] <= 6'h00;
      write_address_data_log_force[7417] <= 6'h00;
      write_address_data_log_force[7418] <= 6'h00;
      write_address_data_log_force[7419] <= 6'h00;
      write_address_data_log_force[7420] <= 6'h00;
      write_address_data_log_force[7421] <= 6'h00;
      write_address_data_log_force[7422] <= 6'h00;
      write_address_data_log_force[7423] <= 6'h00;
      write_address_data_log_force[7424] <= 6'h00;
      write_address_data_log_force[7425] <= 6'h00;
      write_address_data_log_force[7426] <= 6'h00;
      write_address_data_log_force[7427] <= 6'h00;
      write_address_data_log_force[7428] <= 6'h00;
      write_address_data_log_force[7429] <= 6'h00;
      write_address_data_log_force[7430] <= 6'h00;
      write_address_data_log_force[7431] <= 6'h00;
      write_address_data_log_force[7432] <= 6'h00;
      write_address_data_log_force[7433] <= 6'h00;
      write_address_data_log_force[7434] <= 6'h00;
      write_address_data_log_force[7435] <= 6'h00;
      write_address_data_log_force[7436] <= 6'h00;
      write_address_data_log_force[7437] <= 6'h00;
      write_address_data_log_force[7438] <= 6'h00;
      write_address_data_log_force[7439] <= 6'h00;
      write_address_data_log_force[7440] <= 6'h00;
      write_address_data_log_force[7441] <= 6'h00;
      write_address_data_log_force[7442] <= 6'h00;
      write_address_data_log_force[7443] <= 6'h00;
      write_address_data_log_force[7444] <= 6'h00;
      write_address_data_log_force[7445] <= 6'h00;
      write_address_data_log_force[7446] <= 6'h00;
      write_address_data_log_force[7447] <= 6'h00;
      write_address_data_log_force[7448] <= 6'h00;
      write_address_data_log_force[7449] <= 6'h00;
      write_address_data_log_force[7450] <= 6'h00;
      write_address_data_log_force[7451] <= 6'h00;
      write_address_data_log_force[7452] <= 6'h00;
      write_address_data_log_force[7453] <= 6'h00;
      write_address_data_log_force[7454] <= 6'h00;
      write_address_data_log_force[7455] <= 6'h00;
      write_address_data_log_force[7456] <= 6'h00;
      write_address_data_log_force[7457] <= 6'h00;
      write_address_data_log_force[7458] <= 6'h00;
      write_address_data_log_force[7459] <= 6'h00;
      write_address_data_log_force[7460] <= 6'h00;
      write_address_data_log_force[7461] <= 6'h00;
      write_address_data_log_force[7462] <= 6'h00;
      write_address_data_log_force[7463] <= 6'h00;
      write_address_data_log_force[7464] <= 6'h00;
      write_address_data_log_force[7465] <= 6'h00;
      write_address_data_log_force[7466] <= 6'h00;
      write_address_data_log_force[7467] <= 6'h00;
      write_address_data_log_force[7468] <= 6'h00;
      write_address_data_log_force[7469] <= 6'h00;
      write_address_data_log_force[7470] <= 6'h00;
      write_address_data_log_force[7471] <= 6'h00;
      write_address_data_log_force[7472] <= 6'h00;
      write_address_data_log_force[7473] <= 6'h00;
      write_address_data_log_force[7474] <= 6'h00;
      write_address_data_log_force[7475] <= 6'h00;
      write_address_data_log_force[7476] <= 6'h00;
      write_address_data_log_force[7477] <= 6'h00;
      write_address_data_log_force[7478] <= 6'h00;
      write_address_data_log_force[7479] <= 6'h00;
      write_address_data_log_force[7480] <= 6'h00;
      write_address_data_log_force[7481] <= 6'h00;
      write_address_data_log_force[7482] <= 6'h00;
      write_address_data_log_force[7483] <= 6'h00;
      write_address_data_log_force[7484] <= 6'h00;
      write_address_data_log_force[7485] <= 6'h00;
      write_address_data_log_force[7486] <= 6'h00;
      write_address_data_log_force[7487] <= 6'h00;
      write_address_data_log_force[7488] <= 6'h00;
      write_address_data_log_force[7489] <= 6'h00;
      write_address_data_log_force[7490] <= 6'h00;
      write_address_data_log_force[7491] <= 6'h00;
      write_address_data_log_force[7492] <= 6'h00;
      write_address_data_log_force[7493] <= 6'h00;
      write_address_data_log_force[7494] <= 6'h00;
      write_address_data_log_force[7495] <= 6'h00;
      write_address_data_log_force[7496] <= 6'h00;
      write_address_data_log_force[7497] <= 6'h00;
      write_address_data_log_force[7498] <= 6'h00;
      write_address_data_log_force[7499] <= 6'h00;
      write_address_data_log_force[7500] <= 6'h00;
      write_address_data_log_force[7501] <= 6'h00;
      write_address_data_log_force[7502] <= 6'h00;
      write_address_data_log_force[7503] <= 6'h00;
      write_address_data_log_force[7504] <= 6'h00;
      write_address_data_log_force[7505] <= 6'h00;
      write_address_data_log_force[7506] <= 6'h00;
      write_address_data_log_force[7507] <= 6'h00;
      write_address_data_log_force[7508] <= 6'h00;
      write_address_data_log_force[7509] <= 6'h00;
      write_address_data_log_force[7510] <= 6'h00;
      write_address_data_log_force[7511] <= 6'h00;
      write_address_data_log_force[7512] <= 6'h00;
      write_address_data_log_force[7513] <= 6'h00;
      write_address_data_log_force[7514] <= 6'h00;
      write_address_data_log_force[7515] <= 6'h00;
      write_address_data_log_force[7516] <= 6'h00;
      write_address_data_log_force[7517] <= 6'h00;
      write_address_data_log_force[7518] <= 6'h00;
      write_address_data_log_force[7519] <= 6'h00;
      write_address_data_log_force[7520] <= 6'h00;
      write_address_data_log_force[7521] <= 6'h00;
      write_address_data_log_force[7522] <= 6'h00;
      write_address_data_log_force[7523] <= 6'h00;
      write_address_data_log_force[7524] <= 6'h00;
      write_address_data_log_force[7525] <= 6'h00;
      write_address_data_log_force[7526] <= 6'h00;
      write_address_data_log_force[7527] <= 6'h00;
      write_address_data_log_force[7528] <= 6'h00;
      write_address_data_log_force[7529] <= 6'h00;
      write_address_data_log_force[7530] <= 6'h00;
      write_address_data_log_force[7531] <= 6'h00;
      write_address_data_log_force[7532] <= 6'h00;
      write_address_data_log_force[7533] <= 6'h00;
      write_address_data_log_force[7534] <= 6'h00;
      write_address_data_log_force[7535] <= 6'h00;
      write_address_data_log_force[7536] <= 6'h00;
      write_address_data_log_force[7537] <= 6'h00;
      write_address_data_log_force[7538] <= 6'h00;
      write_address_data_log_force[7539] <= 6'h00;
      write_address_data_log_force[7540] <= 6'h00;
      write_address_data_log_force[7541] <= 6'h00;
      write_address_data_log_force[7542] <= 6'h00;
      write_address_data_log_force[7543] <= 6'h00;
      write_address_data_log_force[7544] <= 6'h00;
      write_address_data_log_force[7545] <= 6'h00;
      write_address_data_log_force[7546] <= 6'h00;
      write_address_data_log_force[7547] <= 6'h00;
      write_address_data_log_force[7548] <= 6'h00;
      write_address_data_log_force[7549] <= 6'h00;
      write_address_data_log_force[7550] <= 6'h00;
      write_address_data_log_force[7551] <= 6'h00;
      write_address_data_log_force[7552] <= 6'h00;
      write_address_data_log_force[7553] <= 6'h00;
      write_address_data_log_force[7554] <= 6'h00;
      write_address_data_log_force[7555] <= 6'h00;
      write_address_data_log_force[7556] <= 6'h00;
      write_address_data_log_force[7557] <= 6'h00;
      write_address_data_log_force[7558] <= 6'h00;
      write_address_data_log_force[7559] <= 6'h00;
      write_address_data_log_force[7560] <= 6'h00;
      write_address_data_log_force[7561] <= 6'h00;
      write_address_data_log_force[7562] <= 6'h00;
      write_address_data_log_force[7563] <= 6'h00;
      write_address_data_log_force[7564] <= 6'h00;
      write_address_data_log_force[7565] <= 6'h00;
      write_address_data_log_force[7566] <= 6'h00;
      write_address_data_log_force[7567] <= 6'h00;
      write_address_data_log_force[7568] <= 6'h00;
      write_address_data_log_force[7569] <= 6'h00;
      write_address_data_log_force[7570] <= 6'h00;
      write_address_data_log_force[7571] <= 6'h00;
      write_address_data_log_force[7572] <= 6'h00;
      write_address_data_log_force[7573] <= 6'h00;
      write_address_data_log_force[7574] <= 6'h00;
      write_address_data_log_force[7575] <= 6'h00;
      write_address_data_log_force[7576] <= 6'h00;
      write_address_data_log_force[7577] <= 6'h00;
      write_address_data_log_force[7578] <= 6'h00;
      write_address_data_log_force[7579] <= 6'h00;
      write_address_data_log_force[7580] <= 6'h00;
      write_address_data_log_force[7581] <= 6'h00;
      write_address_data_log_force[7582] <= 6'h00;
      write_address_data_log_force[7583] <= 6'h00;
      write_address_data_log_force[7584] <= 6'h00;
      write_address_data_log_force[7585] <= 6'h00;
      write_address_data_log_force[7586] <= 6'h00;
      write_address_data_log_force[7587] <= 6'h00;
      write_address_data_log_force[7588] <= 6'h00;
      write_address_data_log_force[7589] <= 6'h00;
      write_address_data_log_force[7590] <= 6'h00;
      write_address_data_log_force[7591] <= 6'h00;
      write_address_data_log_force[7592] <= 6'h00;
      write_address_data_log_force[7593] <= 6'h00;
      write_address_data_log_force[7594] <= 6'h00;
      write_address_data_log_force[7595] <= 6'h00;
      write_address_data_log_force[7596] <= 6'h00;
      write_address_data_log_force[7597] <= 6'h00;
      write_address_data_log_force[7598] <= 6'h00;
      write_address_data_log_force[7599] <= 6'h00;
      write_address_data_log_force[7600] <= 6'h00;
      write_address_data_log_force[7601] <= 6'h00;
      write_address_data_log_force[7602] <= 6'h00;
      write_address_data_log_force[7603] <= 6'h00;
      write_address_data_log_force[7604] <= 6'h00;
      write_address_data_log_force[7605] <= 6'h00;
      write_address_data_log_force[7606] <= 6'h00;
      write_address_data_log_force[7607] <= 6'h00;
      write_address_data_log_force[7608] <= 6'h00;
      write_address_data_log_force[7609] <= 6'h00;
      write_address_data_log_force[7610] <= 6'h00;
      write_address_data_log_force[7611] <= 6'h00;
      write_address_data_log_force[7612] <= 6'h00;
      write_address_data_log_force[7613] <= 6'h00;
      write_address_data_log_force[7614] <= 6'h00;
      write_address_data_log_force[7615] <= 6'h00;
      write_address_data_log_force[7616] <= 6'h00;
      write_address_data_log_force[7617] <= 6'h00;
      write_address_data_log_force[7618] <= 6'h00;
      write_address_data_log_force[7619] <= 6'h00;
      write_address_data_log_force[7620] <= 6'h00;
      write_address_data_log_force[7621] <= 6'h00;
      write_address_data_log_force[7622] <= 6'h00;
      write_address_data_log_force[7623] <= 6'h00;
      write_address_data_log_force[7624] <= 6'h00;
      write_address_data_log_force[7625] <= 6'h00;
      write_address_data_log_force[7626] <= 6'h00;
      write_address_data_log_force[7627] <= 6'h00;
      write_address_data_log_force[7628] <= 6'h00;
      write_address_data_log_force[7629] <= 6'h00;
      write_address_data_log_force[7630] <= 6'h00;
      write_address_data_log_force[7631] <= 6'h00;
      write_address_data_log_force[7632] <= 6'h00;
      write_address_data_log_force[7633] <= 6'h00;
      write_address_data_log_force[7634] <= 6'h00;
      write_address_data_log_force[7635] <= 6'h00;
      write_address_data_log_force[7636] <= 6'h00;
      write_address_data_log_force[7637] <= 6'h00;
      write_address_data_log_force[7638] <= 6'h00;
      write_address_data_log_force[7639] <= 6'h00;
      write_address_data_log_force[7640] <= 6'h00;
      write_address_data_log_force[7641] <= 6'h00;
      write_address_data_log_force[7642] <= 6'h00;
      write_address_data_log_force[7643] <= 6'h00;
      write_address_data_log_force[7644] <= 6'h00;
      write_address_data_log_force[7645] <= 6'h00;
      write_address_data_log_force[7646] <= 6'h00;
      write_address_data_log_force[7647] <= 6'h00;
      write_address_data_log_force[7648] <= 6'h00;
      write_address_data_log_force[7649] <= 6'h00;
      write_address_data_log_force[7650] <= 6'h00;
      write_address_data_log_force[7651] <= 6'h00;
      write_address_data_log_force[7652] <= 6'h00;
      write_address_data_log_force[7653] <= 6'h00;
      write_address_data_log_force[7654] <= 6'h00;
      write_address_data_log_force[7655] <= 6'h00;
      write_address_data_log_force[7656] <= 6'h00;
      write_address_data_log_force[7657] <= 6'h00;
      write_address_data_log_force[7658] <= 6'h00;
      write_address_data_log_force[7659] <= 6'h00;
      write_address_data_log_force[7660] <= 6'h00;
      write_address_data_log_force[7661] <= 6'h00;
      write_address_data_log_force[7662] <= 6'h00;
      write_address_data_log_force[7663] <= 6'h00;
      write_address_data_log_force[7664] <= 6'h00;
      write_address_data_log_force[7665] <= 6'h00;
      write_address_data_log_force[7666] <= 6'h00;
      write_address_data_log_force[7667] <= 6'h00;
      write_address_data_log_force[7668] <= 6'h00;
      write_address_data_log_force[7669] <= 6'h00;
      write_address_data_log_force[7670] <= 6'h00;
      write_address_data_log_force[7671] <= 6'h00;
      write_address_data_log_force[7672] <= 6'h00;
      write_address_data_log_force[7673] <= 6'h00;
      write_address_data_log_force[7674] <= 6'h00;
      write_address_data_log_force[7675] <= 6'h00;
      write_address_data_log_force[7676] <= 6'h00;
      write_address_data_log_force[7677] <= 6'h00;
      write_address_data_log_force[7678] <= 6'h00;
      write_address_data_log_force[7679] <= 6'h00;
      write_address_data_log_force[7680] <= 6'h00;
      write_address_data_log_force[7681] <= 6'h00;
      write_address_data_log_force[7682] <= 6'h00;
      write_address_data_log_force[7683] <= 6'h00;
      write_address_data_log_force[7684] <= 6'h00;
      write_address_data_log_force[7685] <= 6'h00;
      write_address_data_log_force[7686] <= 6'h00;
      write_address_data_log_force[7687] <= 6'h00;
      write_address_data_log_force[7688] <= 6'h00;
      write_address_data_log_force[7689] <= 6'h00;
      write_address_data_log_force[7690] <= 6'h00;
      write_address_data_log_force[7691] <= 6'h00;
      write_address_data_log_force[7692] <= 6'h00;
      write_address_data_log_force[7693] <= 6'h00;
      write_address_data_log_force[7694] <= 6'h00;
      write_address_data_log_force[7695] <= 6'h00;
      write_address_data_log_force[7696] <= 6'h00;
      write_address_data_log_force[7697] <= 6'h00;
      write_address_data_log_force[7698] <= 6'h00;
      write_address_data_log_force[7699] <= 6'h00;
      write_address_data_log_force[7700] <= 6'h00;
      write_address_data_log_force[7701] <= 6'h00;
      write_address_data_log_force[7702] <= 6'h00;
      write_address_data_log_force[7703] <= 6'h00;
      write_address_data_log_force[7704] <= 6'h00;
      write_address_data_log_force[7705] <= 6'h00;
      write_address_data_log_force[7706] <= 6'h00;
      write_address_data_log_force[7707] <= 6'h00;
      write_address_data_log_force[7708] <= 6'h00;
      write_address_data_log_force[7709] <= 6'h00;
      write_address_data_log_force[7710] <= 6'h00;
      write_address_data_log_force[7711] <= 6'h00;
      write_address_data_log_force[7712] <= 6'h00;
      write_address_data_log_force[7713] <= 6'h00;
      write_address_data_log_force[7714] <= 6'h00;
      write_address_data_log_force[7715] <= 6'h00;
      write_address_data_log_force[7716] <= 6'h00;
      write_address_data_log_force[7717] <= 6'h00;
      write_address_data_log_force[7718] <= 6'h00;
      write_address_data_log_force[7719] <= 6'h00;
      write_address_data_log_force[7720] <= 6'h00;
      write_address_data_log_force[7721] <= 6'h00;
      write_address_data_log_force[7722] <= 6'h00;
      write_address_data_log_force[7723] <= 6'h00;
      write_address_data_log_force[7724] <= 6'h00;
      write_address_data_log_force[7725] <= 6'h00;
      write_address_data_log_force[7726] <= 6'h00;
      write_address_data_log_force[7727] <= 6'h00;
      write_address_data_log_force[7728] <= 6'h00;
      write_address_data_log_force[7729] <= 6'h00;
      write_address_data_log_force[7730] <= 6'h00;
      write_address_data_log_force[7731] <= 6'h00;
      write_address_data_log_force[7732] <= 6'h00;
      write_address_data_log_force[7733] <= 6'h00;
      write_address_data_log_force[7734] <= 6'h00;
      write_address_data_log_force[7735] <= 6'h00;
      write_address_data_log_force[7736] <= 6'h00;
      write_address_data_log_force[7737] <= 6'h00;
      write_address_data_log_force[7738] <= 6'h00;
      write_address_data_log_force[7739] <= 6'h00;
      write_address_data_log_force[7740] <= 6'h00;
      write_address_data_log_force[7741] <= 6'h00;
      write_address_data_log_force[7742] <= 6'h00;
      write_address_data_log_force[7743] <= 6'h00;
      write_address_data_log_force[7744] <= 6'h00;
      write_address_data_log_force[7745] <= 6'h00;
      write_address_data_log_force[7746] <= 6'h00;
      write_address_data_log_force[7747] <= 6'h00;
      write_address_data_log_force[7748] <= 6'h00;
      write_address_data_log_force[7749] <= 6'h00;
      write_address_data_log_force[7750] <= 6'h00;
      write_address_data_log_force[7751] <= 6'h00;
      write_address_data_log_force[7752] <= 6'h00;
      write_address_data_log_force[7753] <= 6'h00;
      write_address_data_log_force[7754] <= 6'h00;
      write_address_data_log_force[7755] <= 6'h00;
      write_address_data_log_force[7756] <= 6'h00;
      write_address_data_log_force[7757] <= 6'h00;
      write_address_data_log_force[7758] <= 6'h00;
      write_address_data_log_force[7759] <= 6'h00;
      write_address_data_log_force[7760] <= 6'h00;
      write_address_data_log_force[7761] <= 6'h00;
      write_address_data_log_force[7762] <= 6'h00;
      write_address_data_log_force[7763] <= 6'h00;
      write_address_data_log_force[7764] <= 6'h00;
      write_address_data_log_force[7765] <= 6'h00;
      write_address_data_log_force[7766] <= 6'h00;
      write_address_data_log_force[7767] <= 6'h00;
      write_address_data_log_force[7768] <= 6'h00;
      write_address_data_log_force[7769] <= 6'h00;
      write_address_data_log_force[7770] <= 6'h00;
      write_address_data_log_force[7771] <= 6'h00;
      write_address_data_log_force[7772] <= 6'h00;
      write_address_data_log_force[7773] <= 6'h00;
      write_address_data_log_force[7774] <= 6'h00;
      write_address_data_log_force[7775] <= 6'h00;
      write_address_data_log_force[7776] <= 6'h00;
      write_address_data_log_force[7777] <= 6'h00;
      write_address_data_log_force[7778] <= 6'h00;
      write_address_data_log_force[7779] <= 6'h00;
      write_address_data_log_force[7780] <= 6'h00;
      write_address_data_log_force[7781] <= 6'h00;
      write_address_data_log_force[7782] <= 6'h00;
      write_address_data_log_force[7783] <= 6'h00;
      write_address_data_log_force[7784] <= 6'h00;
      write_address_data_log_force[7785] <= 6'h00;
      write_address_data_log_force[7786] <= 6'h00;
      write_address_data_log_force[7787] <= 6'h00;
      write_address_data_log_force[7788] <= 6'h00;
      write_address_data_log_force[7789] <= 6'h00;
      write_address_data_log_force[7790] <= 6'h00;
      write_address_data_log_force[7791] <= 6'h00;
      write_address_data_log_force[7792] <= 6'h00;
      write_address_data_log_force[7793] <= 6'h00;
      write_address_data_log_force[7794] <= 6'h00;
      write_address_data_log_force[7795] <= 6'h00;
      write_address_data_log_force[7796] <= 6'h00;
      write_address_data_log_force[7797] <= 6'h00;
      write_address_data_log_force[7798] <= 6'h00;
      write_address_data_log_force[7799] <= 6'h00;
      write_address_data_log_force[7800] <= 6'h00;
      write_address_data_log_force[7801] <= 6'h00;
      write_address_data_log_force[7802] <= 6'h00;
      write_address_data_log_force[7803] <= 6'h00;
      write_address_data_log_force[7804] <= 6'h00;
      write_address_data_log_force[7805] <= 6'h00;
      write_address_data_log_force[7806] <= 6'h00;
      write_address_data_log_force[7807] <= 6'h00;
      write_address_data_log_force[7808] <= 6'h00;
      write_address_data_log_force[7809] <= 6'h00;
      write_address_data_log_force[7810] <= 6'h00;
      write_address_data_log_force[7811] <= 6'h00;
      write_address_data_log_force[7812] <= 6'h00;
      write_address_data_log_force[7813] <= 6'h00;
      write_address_data_log_force[7814] <= 6'h00;
      write_address_data_log_force[7815] <= 6'h00;
      write_address_data_log_force[7816] <= 6'h00;
      write_address_data_log_force[7817] <= 6'h00;
      write_address_data_log_force[7818] <= 6'h00;
      write_address_data_log_force[7819] <= 6'h00;
      write_address_data_log_force[7820] <= 6'h00;
      write_address_data_log_force[7821] <= 6'h00;
      write_address_data_log_force[7822] <= 6'h00;
      write_address_data_log_force[7823] <= 6'h00;
      write_address_data_log_force[7824] <= 6'h00;
      write_address_data_log_force[7825] <= 6'h00;
      write_address_data_log_force[7826] <= 6'h00;
      write_address_data_log_force[7827] <= 6'h00;
      write_address_data_log_force[7828] <= 6'h00;
      write_address_data_log_force[7829] <= 6'h00;
      write_address_data_log_force[7830] <= 6'h00;
      write_address_data_log_force[7831] <= 6'h00;
      write_address_data_log_force[7832] <= 6'h00;
      write_address_data_log_force[7833] <= 6'h00;
      write_address_data_log_force[7834] <= 6'h00;
      write_address_data_log_force[7835] <= 6'h00;
      write_address_data_log_force[7836] <= 6'h00;
      write_address_data_log_force[7837] <= 6'h00;
      write_address_data_log_force[7838] <= 6'h00;
      write_address_data_log_force[7839] <= 6'h00;
      write_address_data_log_force[7840] <= 6'h00;
      write_address_data_log_force[7841] <= 6'h00;
      write_address_data_log_force[7842] <= 6'h00;
      write_address_data_log_force[7843] <= 6'h00;
      write_address_data_log_force[7844] <= 6'h00;
      write_address_data_log_force[7845] <= 6'h00;
      write_address_data_log_force[7846] <= 6'h00;
      write_address_data_log_force[7847] <= 6'h00;
      write_address_data_log_force[7848] <= 6'h00;
      write_address_data_log_force[7849] <= 6'h00;
      write_address_data_log_force[7850] <= 6'h00;
      write_address_data_log_force[7851] <= 6'h00;
      write_address_data_log_force[7852] <= 6'h00;
      write_address_data_log_force[7853] <= 6'h00;
      write_address_data_log_force[7854] <= 6'h00;
      write_address_data_log_force[7855] <= 6'h00;
      write_address_data_log_force[7856] <= 6'h00;
      write_address_data_log_force[7857] <= 6'h00;
      write_address_data_log_force[7858] <= 6'h00;
      write_address_data_log_force[7859] <= 6'h00;
      write_address_data_log_force[7860] <= 6'h00;
      write_address_data_log_force[7861] <= 6'h00;
      write_address_data_log_force[7862] <= 6'h00;
      write_address_data_log_force[7863] <= 6'h00;
      write_address_data_log_force[7864] <= 6'h00;
      write_address_data_log_force[7865] <= 6'h00;
      write_address_data_log_force[7866] <= 6'h00;
      write_address_data_log_force[7867] <= 6'h00;
      write_address_data_log_force[7868] <= 6'h00;
      write_address_data_log_force[7869] <= 6'h00;
      write_address_data_log_force[7870] <= 6'h00;
      write_address_data_log_force[7871] <= 6'h00;
      write_address_data_log_force[7872] <= 6'h00;
      write_address_data_log_force[7873] <= 6'h00;
      write_address_data_log_force[7874] <= 6'h00;
      write_address_data_log_force[7875] <= 6'h00;
      write_address_data_log_force[7876] <= 6'h00;
      write_address_data_log_force[7877] <= 6'h00;
      write_address_data_log_force[7878] <= 6'h00;
      write_address_data_log_force[7879] <= 6'h00;
      write_address_data_log_force[7880] <= 6'h00;
      write_address_data_log_force[7881] <= 6'h00;
      write_address_data_log_force[7882] <= 6'h00;
      write_address_data_log_force[7883] <= 6'h00;
      write_address_data_log_force[7884] <= 6'h00;
      write_address_data_log_force[7885] <= 6'h00;
      write_address_data_log_force[7886] <= 6'h00;
      write_address_data_log_force[7887] <= 6'h00;
      write_address_data_log_force[7888] <= 6'h00;
      write_address_data_log_force[7889] <= 6'h00;
      write_address_data_log_force[7890] <= 6'h00;
      write_address_data_log_force[7891] <= 6'h00;
      write_address_data_log_force[7892] <= 6'h00;
      write_address_data_log_force[7893] <= 6'h00;
      write_address_data_log_force[7894] <= 6'h00;
      write_address_data_log_force[7895] <= 6'h00;
      write_address_data_log_force[7896] <= 6'h00;
      write_address_data_log_force[7897] <= 6'h00;
      write_address_data_log_force[7898] <= 6'h00;
      write_address_data_log_force[7899] <= 6'h00;
      write_address_data_log_force[7900] <= 6'h00;
      write_address_data_log_force[7901] <= 6'h00;
      write_address_data_log_force[7902] <= 6'h00;
      write_address_data_log_force[7903] <= 6'h00;
      write_address_data_log_force[7904] <= 6'h00;
      write_address_data_log_force[7905] <= 6'h00;
      write_address_data_log_force[7906] <= 6'h00;
      write_address_data_log_force[7907] <= 6'h00;
      write_address_data_log_force[7908] <= 6'h00;
      write_address_data_log_force[7909] <= 6'h00;
      write_address_data_log_force[7910] <= 6'h00;
      write_address_data_log_force[7911] <= 6'h00;
      write_address_data_log_force[7912] <= 6'h00;
      write_address_data_log_force[7913] <= 6'h00;
      write_address_data_log_force[7914] <= 6'h00;
      write_address_data_log_force[7915] <= 6'h00;
      write_address_data_log_force[7916] <= 6'h00;
      write_address_data_log_force[7917] <= 6'h00;
      write_address_data_log_force[7918] <= 6'h00;
      write_address_data_log_force[7919] <= 6'h00;
      write_address_data_log_force[7920] <= 6'h00;
      write_address_data_log_force[7921] <= 6'h00;
      write_address_data_log_force[7922] <= 6'h00;
      write_address_data_log_force[7923] <= 6'h00;
      write_address_data_log_force[7924] <= 6'h00;
      write_address_data_log_force[7925] <= 6'h00;
      write_address_data_log_force[7926] <= 6'h00;
      write_address_data_log_force[7927] <= 6'h00;
      write_address_data_log_force[7928] <= 6'h00;
      write_address_data_log_force[7929] <= 6'h00;
      write_address_data_log_force[7930] <= 6'h00;
      write_address_data_log_force[7931] <= 6'h00;
      write_address_data_log_force[7932] <= 6'h00;
      write_address_data_log_force[7933] <= 6'h00;
      write_address_data_log_force[7934] <= 6'h00;
      write_address_data_log_force[7935] <= 6'h00;
      write_address_data_log_force[7936] <= 6'h00;
      write_address_data_log_force[7937] <= 6'h00;
      write_address_data_log_force[7938] <= 6'h00;
      write_address_data_log_force[7939] <= 6'h00;
      write_address_data_log_force[7940] <= 6'h00;
      write_address_data_log_force[7941] <= 6'h00;
      write_address_data_log_force[7942] <= 6'h00;
      write_address_data_log_force[7943] <= 6'h00;
      write_address_data_log_force[7944] <= 6'h00;
      write_address_data_log_force[7945] <= 6'h00;
      write_address_data_log_force[7946] <= 6'h00;
      write_address_data_log_force[7947] <= 6'h00;
      write_address_data_log_force[7948] <= 6'h00;
      write_address_data_log_force[7949] <= 6'h00;
      write_address_data_log_force[7950] <= 6'h00;
      write_address_data_log_force[7951] <= 6'h00;
      write_address_data_log_force[7952] <= 6'h00;
      write_address_data_log_force[7953] <= 6'h00;
      write_address_data_log_force[7954] <= 6'h00;
      write_address_data_log_force[7955] <= 6'h00;
      write_address_data_log_force[7956] <= 6'h00;
      write_address_data_log_force[7957] <= 6'h00;
      write_address_data_log_force[7958] <= 6'h00;
      write_address_data_log_force[7959] <= 6'h00;
      write_address_data_log_force[7960] <= 6'h00;
      write_address_data_log_force[7961] <= 6'h00;
      write_address_data_log_force[7962] <= 6'h00;
      write_address_data_log_force[7963] <= 6'h00;
      write_address_data_log_force[7964] <= 6'h00;
      write_address_data_log_force[7965] <= 6'h00;
      write_address_data_log_force[7966] <= 6'h00;
      write_address_data_log_force[7967] <= 6'h00;
      write_address_data_log_force[7968] <= 6'h00;
      write_address_data_log_force[7969] <= 6'h00;
      write_address_data_log_force[7970] <= 6'h00;
      write_address_data_log_force[7971] <= 6'h00;
      write_address_data_log_force[7972] <= 6'h00;
      write_address_data_log_force[7973] <= 6'h00;
      write_address_data_log_force[7974] <= 6'h00;
      write_address_data_log_force[7975] <= 6'h00;
      write_address_data_log_force[7976] <= 6'h00;
      write_address_data_log_force[7977] <= 6'h00;
      write_address_data_log_force[7978] <= 6'h00;
      write_address_data_log_force[7979] <= 6'h00;
      write_address_data_log_force[7980] <= 6'h00;
      write_address_data_log_force[7981] <= 6'h00;
      write_address_data_log_force[7982] <= 6'h00;
      write_address_data_log_force[7983] <= 6'h00;
      write_address_data_log_force[7984] <= 6'h00;
      write_address_data_log_force[7985] <= 6'h00;
      write_address_data_log_force[7986] <= 6'h00;
      write_address_data_log_force[7987] <= 6'h00;
      write_address_data_log_force[7988] <= 6'h00;
      write_address_data_log_force[7989] <= 6'h00;
      write_address_data_log_force[7990] <= 6'h00;
      write_address_data_log_force[7991] <= 6'h00;
      write_address_data_log_force[7992] <= 6'h00;
      write_address_data_log_force[7993] <= 6'h00;
      write_address_data_log_force[7994] <= 6'h00;
      write_address_data_log_force[7995] <= 6'h00;
      write_address_data_log_force[7996] <= 6'h00;
      write_address_data_log_force[7997] <= 6'h00;
      write_address_data_log_force[7998] <= 6'h00;
      write_address_data_log_force[7999] <= 6'h00;
      write_address_data_log_force[8000] <= 6'h00;
      write_address_data_log_force[8001] <= 6'h00;
      write_address_data_log_force[8002] <= 6'h00;
      write_address_data_log_force[8003] <= 6'h00;
      write_address_data_log_force[8004] <= 6'h00;
      write_address_data_log_force[8005] <= 6'h00;
      write_address_data_log_force[8006] <= 6'h00;
      write_address_data_log_force[8007] <= 6'h00;
      write_address_data_log_force[8008] <= 6'h00;
      write_address_data_log_force[8009] <= 6'h00;
      write_address_data_log_force[8010] <= 6'h00;
      write_address_data_log_force[8011] <= 6'h00;
      write_address_data_log_force[8012] <= 6'h00;
      write_address_data_log_force[8013] <= 6'h00;
      write_address_data_log_force[8014] <= 6'h00;
      write_address_data_log_force[8015] <= 6'h00;
      write_address_data_log_force[8016] <= 6'h00;
      write_address_data_log_force[8017] <= 6'h00;
      write_address_data_log_force[8018] <= 6'h00;
      write_address_data_log_force[8019] <= 6'h00;
      write_address_data_log_force[8020] <= 6'h00;
      write_address_data_log_force[8021] <= 6'h00;
      write_address_data_log_force[8022] <= 6'h00;
      write_address_data_log_force[8023] <= 6'h00;
      write_address_data_log_force[8024] <= 6'h00;
      write_address_data_log_force[8025] <= 6'h00;
      write_address_data_log_force[8026] <= 6'h00;
      write_address_data_log_force[8027] <= 6'h00;
      write_address_data_log_force[8028] <= 6'h00;
      write_address_data_log_force[8029] <= 6'h00;
      write_address_data_log_force[8030] <= 6'h00;
      write_address_data_log_force[8031] <= 6'h00;
      write_address_data_log_force[8032] <= 6'h00;
      write_address_data_log_force[8033] <= 6'h00;
      write_address_data_log_force[8034] <= 6'h00;
      write_address_data_log_force[8035] <= 6'h00;
      write_address_data_log_force[8036] <= 6'h00;
      write_address_data_log_force[8037] <= 6'h00;
      write_address_data_log_force[8038] <= 6'h00;
      write_address_data_log_force[8039] <= 6'h00;
      write_address_data_log_force[8040] <= 6'h00;
      write_address_data_log_force[8041] <= 6'h00;
      write_address_data_log_force[8042] <= 6'h00;
      write_address_data_log_force[8043] <= 6'h00;
      write_address_data_log_force[8044] <= 6'h00;
      write_address_data_log_force[8045] <= 6'h00;
      write_address_data_log_force[8046] <= 6'h00;
      write_address_data_log_force[8047] <= 6'h00;
      write_address_data_log_force[8048] <= 6'h00;
      write_address_data_log_force[8049] <= 6'h00;
      write_address_data_log_force[8050] <= 6'h00;
      write_address_data_log_force[8051] <= 6'h00;
      write_address_data_log_force[8052] <= 6'h00;
      write_address_data_log_force[8053] <= 6'h00;
      write_address_data_log_force[8054] <= 6'h00;
      write_address_data_log_force[8055] <= 6'h00;
      write_address_data_log_force[8056] <= 6'h00;
      write_address_data_log_force[8057] <= 6'h00;
      write_address_data_log_force[8058] <= 6'h00;
      write_address_data_log_force[8059] <= 6'h00;
      write_address_data_log_force[8060] <= 6'h00;
      write_address_data_log_force[8061] <= 6'h00;
      write_address_data_log_force[8062] <= 6'h00;
      write_address_data_log_force[8063] <= 6'h00;
      write_address_data_log_force[8064] <= 6'h00;
      write_address_data_log_force[8065] <= 6'h00;
      write_address_data_log_force[8066] <= 6'h00;
      write_address_data_log_force[8067] <= 6'h00;
      write_address_data_log_force[8068] <= 6'h00;
      write_address_data_log_force[8069] <= 6'h00;
      write_address_data_log_force[8070] <= 6'h00;
      write_address_data_log_force[8071] <= 6'h00;
      write_address_data_log_force[8072] <= 6'h00;
      write_address_data_log_force[8073] <= 6'h00;
      write_address_data_log_force[8074] <= 6'h00;
      write_address_data_log_force[8075] <= 6'h00;
      write_address_data_log_force[8076] <= 6'h00;
      write_address_data_log_force[8077] <= 6'h00;
      write_address_data_log_force[8078] <= 6'h00;
      write_address_data_log_force[8079] <= 6'h00;
      write_address_data_log_force[8080] <= 6'h00;
      write_address_data_log_force[8081] <= 6'h00;
      write_address_data_log_force[8082] <= 6'h00;
      write_address_data_log_force[8083] <= 6'h00;
      write_address_data_log_force[8084] <= 6'h00;
      write_address_data_log_force[8085] <= 6'h00;
      write_address_data_log_force[8086] <= 6'h00;
      write_address_data_log_force[8087] <= 6'h00;
      write_address_data_log_force[8088] <= 6'h00;
      write_address_data_log_force[8089] <= 6'h00;
      write_address_data_log_force[8090] <= 6'h00;
      write_address_data_log_force[8091] <= 6'h00;
      write_address_data_log_force[8092] <= 6'h00;
      write_address_data_log_force[8093] <= 6'h00;
      write_address_data_log_force[8094] <= 6'h00;
      write_address_data_log_force[8095] <= 6'h00;
      write_address_data_log_force[8096] <= 6'h00;
      write_address_data_log_force[8097] <= 6'h00;
      write_address_data_log_force[8098] <= 6'h00;
      write_address_data_log_force[8099] <= 6'h00;
      write_address_data_log_force[8100] <= 6'h00;
      write_address_data_log_force[8101] <= 6'h00;
      write_address_data_log_force[8102] <= 6'h00;
      write_address_data_log_force[8103] <= 6'h00;
      write_address_data_log_force[8104] <= 6'h00;
      write_address_data_log_force[8105] <= 6'h00;
      write_address_data_log_force[8106] <= 6'h00;
      write_address_data_log_force[8107] <= 6'h00;
      write_address_data_log_force[8108] <= 6'h00;
      write_address_data_log_force[8109] <= 6'h00;
      write_address_data_log_force[8110] <= 6'h00;
      write_address_data_log_force[8111] <= 6'h00;
      write_address_data_log_force[8112] <= 6'h00;
      write_address_data_log_force[8113] <= 6'h00;
      write_address_data_log_force[8114] <= 6'h00;
      write_address_data_log_force[8115] <= 6'h00;
      write_address_data_log_force[8116] <= 6'h00;
      write_address_data_log_force[8117] <= 6'h00;
      write_address_data_log_force[8118] <= 6'h00;
      write_address_data_log_force[8119] <= 6'h00;
      write_address_data_log_force[8120] <= 6'h00;
      write_address_data_log_force[8121] <= 6'h00;
      write_address_data_log_force[8122] <= 6'h00;
      write_address_data_log_force[8123] <= 6'h00;
      write_address_data_log_force[8124] <= 6'h00;
      write_address_data_log_force[8125] <= 6'h00;
      write_address_data_log_force[8126] <= 6'h00;
      write_address_data_log_force[8127] <= 6'h00;
      write_address_data_log_force[8128] <= 6'h00;
      write_address_data_log_force[8129] <= 6'h00;
      write_address_data_log_force[8130] <= 6'h00;
      write_address_data_log_force[8131] <= 6'h00;
      write_address_data_log_force[8132] <= 6'h00;
      write_address_data_log_force[8133] <= 6'h00;
      write_address_data_log_force[8134] <= 6'h00;
      write_address_data_log_force[8135] <= 6'h00;
      write_address_data_log_force[8136] <= 6'h00;
      write_address_data_log_force[8137] <= 6'h00;
      write_address_data_log_force[8138] <= 6'h00;
      write_address_data_log_force[8139] <= 6'h00;
      write_address_data_log_force[8140] <= 6'h00;
      write_address_data_log_force[8141] <= 6'h00;
      write_address_data_log_force[8142] <= 6'h00;
      write_address_data_log_force[8143] <= 6'h00;
      write_address_data_log_force[8144] <= 6'h00;
      write_address_data_log_force[8145] <= 6'h00;
      write_address_data_log_force[8146] <= 6'h00;
      write_address_data_log_force[8147] <= 6'h00;
      write_address_data_log_force[8148] <= 6'h00;
      write_address_data_log_force[8149] <= 6'h00;
      write_address_data_log_force[8150] <= 6'h00;
      write_address_data_log_force[8151] <= 6'h00;
      write_address_data_log_force[8152] <= 6'h00;
      write_address_data_log_force[8153] <= 6'h00;
      write_address_data_log_force[8154] <= 6'h00;
      write_address_data_log_force[8155] <= 6'h00;
      write_address_data_log_force[8156] <= 6'h00;
      write_address_data_log_force[8157] <= 6'h00;
      write_address_data_log_force[8158] <= 6'h00;
      write_address_data_log_force[8159] <= 6'h00;
      write_address_data_log_force[8160] <= 6'h00;
      write_address_data_log_force[8161] <= 6'h00;
      write_address_data_log_force[8162] <= 6'h00;
      write_address_data_log_force[8163] <= 6'h00;
      write_address_data_log_force[8164] <= 6'h00;
      write_address_data_log_force[8165] <= 6'h00;
      write_address_data_log_force[8166] <= 6'h00;
      write_address_data_log_force[8167] <= 6'h00;
      write_address_data_log_force[8168] <= 6'h00;
      write_address_data_log_force[8169] <= 6'h00;
      write_address_data_log_force[8170] <= 6'h00;
      write_address_data_log_force[8171] <= 6'h00;
      write_address_data_log_force[8172] <= 6'h00;
      write_address_data_log_force[8173] <= 6'h00;
      write_address_data_log_force[8174] <= 6'h00;
      write_address_data_log_force[8175] <= 6'h00;
      write_address_data_log_force[8176] <= 6'h00;
      write_address_data_log_force[8177] <= 6'h00;
      write_address_data_log_force[8178] <= 6'h00;
      write_address_data_log_force[8179] <= 6'h00;
      write_address_data_log_force[8180] <= 6'h00;
      write_address_data_log_force[8181] <= 6'h00;
      write_address_data_log_force[8182] <= 6'h00;
      write_address_data_log_force[8183] <= 6'h00;
      write_address_data_log_force[8184] <= 6'h00;
      write_address_data_log_force[8185] <= 6'h00;
      write_address_data_log_force[8186] <= 6'h00;
      write_address_data_log_force[8187] <= 6'h00;
      write_address_data_log_force[8188] <= 6'h00;
      write_address_data_log_force[8189] <= 6'h00;
      write_address_data_log_force[8190] <= 6'h00;
      write_address_data_log_force[8191] <= 6'h00;
      write_address_data_log_force[8192] <= 6'h00;
      write_address_data_log_force[8193] <= 6'h00;
      write_address_data_log_force[8194] <= 6'h00;
      write_address_data_log_force[8195] <= 6'h00;
      write_address_data_log_force[8196] <= 6'h00;
      write_address_data_log_force[8197] <= 6'h00;
      write_address_data_log_force[8198] <= 6'h00;
      write_address_data_log_force[8199] <= 6'h00;
      write_address_data_log_force[8200] <= 6'h00;
      write_address_data_log_force[8201] <= 6'h00;
      write_address_data_log_force[8202] <= 6'h00;
      write_address_data_log_force[8203] <= 6'h00;
      write_address_data_log_force[8204] <= 6'h00;
      write_address_data_log_force[8205] <= 6'h00;
      write_address_data_log_force[8206] <= 6'h00;
      write_address_data_log_force[8207] <= 6'h00;
      write_address_data_log_force[8208] <= 6'h00;
      write_address_data_log_force[8209] <= 6'h00;
      write_address_data_log_force[8210] <= 6'h00;
      write_address_data_log_force[8211] <= 6'h00;
      write_address_data_log_force[8212] <= 6'h00;
      write_address_data_log_force[8213] <= 6'h00;
      write_address_data_log_force[8214] <= 6'h00;
      write_address_data_log_force[8215] <= 6'h00;
      write_address_data_log_force[8216] <= 6'h00;
      write_address_data_log_force[8217] <= 6'h00;
      write_address_data_log_force[8218] <= 6'h00;
      write_address_data_log_force[8219] <= 6'h00;
      write_address_data_log_force[8220] <= 6'h00;
      write_address_data_log_force[8221] <= 6'h00;
      write_address_data_log_force[8222] <= 6'h00;
      write_address_data_log_force[8223] <= 6'h00;
      write_address_data_log_force[8224] <= 6'h00;
      write_address_data_log_force[8225] <= 6'h00;
      write_address_data_log_force[8226] <= 6'h00;
      write_address_data_log_force[8227] <= 6'h00;
      write_address_data_log_force[8228] <= 6'h00;
      write_address_data_log_force[8229] <= 6'h00;
      write_address_data_log_force[8230] <= 6'h00;
      write_address_data_log_force[8231] <= 6'h00;
      write_address_data_log_force[8232] <= 6'h00;
      write_address_data_log_force[8233] <= 6'h00;
      write_address_data_log_force[8234] <= 6'h00;
      write_address_data_log_force[8235] <= 6'h00;
      write_address_data_log_force[8236] <= 6'h00;
      write_address_data_log_force[8237] <= 6'h00;
      write_address_data_log_force[8238] <= 6'h00;
      write_address_data_log_force[8239] <= 6'h00;
      write_address_data_log_force[8240] <= 6'h00;
      write_address_data_log_force[8241] <= 6'h00;
      write_address_data_log_force[8242] <= 6'h00;
      write_address_data_log_force[8243] <= 6'h00;
      write_address_data_log_force[8244] <= 6'h00;
      write_address_data_log_force[8245] <= 6'h00;
      write_address_data_log_force[8246] <= 6'h00;
      write_address_data_log_force[8247] <= 6'h00;
      write_address_data_log_force[8248] <= 6'h00;
      write_address_data_log_force[8249] <= 6'h00;
      write_address_data_log_force[8250] <= 6'h00;
      write_address_data_log_force[8251] <= 6'h00;
      write_address_data_log_force[8252] <= 6'h00;
      write_address_data_log_force[8253] <= 6'h00;
      write_address_data_log_force[8254] <= 6'h00;
      write_address_data_log_force[8255] <= 6'h00;
      write_address_data_log_force[8256] <= 6'h00;
      write_address_data_log_force[8257] <= 6'h00;
      write_address_data_log_force[8258] <= 6'h00;
      write_address_data_log_force[8259] <= 6'h00;
      write_address_data_log_force[8260] <= 6'h00;
      write_address_data_log_force[8261] <= 6'h00;
      write_address_data_log_force[8262] <= 6'h00;
      write_address_data_log_force[8263] <= 6'h00;
      write_address_data_log_force[8264] <= 6'h00;
      write_address_data_log_force[8265] <= 6'h00;
      write_address_data_log_force[8266] <= 6'h00;
      write_address_data_log_force[8267] <= 6'h00;
      write_address_data_log_force[8268] <= 6'h00;
      write_address_data_log_force[8269] <= 6'h00;
      write_address_data_log_force[8270] <= 6'h00;
      write_address_data_log_force[8271] <= 6'h00;
      write_address_data_log_force[8272] <= 6'h00;
      write_address_data_log_force[8273] <= 6'h00;
      write_address_data_log_force[8274] <= 6'h00;
      write_address_data_log_force[8275] <= 6'h00;
      write_address_data_log_force[8276] <= 6'h00;
      write_address_data_log_force[8277] <= 6'h00;
      write_address_data_log_force[8278] <= 6'h00;
      write_address_data_log_force[8279] <= 6'h00;
      write_address_data_log_force[8280] <= 6'h00;
      write_address_data_log_force[8281] <= 6'h00;
      write_address_data_log_force[8282] <= 6'h00;
      write_address_data_log_force[8283] <= 6'h00;
      write_address_data_log_force[8284] <= 6'h00;
      write_address_data_log_force[8285] <= 6'h00;
      write_address_data_log_force[8286] <= 6'h00;
      write_address_data_log_force[8287] <= 6'h00;
      write_address_data_log_force[8288] <= 6'h00;
      write_address_data_log_force[8289] <= 6'h00;
      write_address_data_log_force[8290] <= 6'h00;
      write_address_data_log_force[8291] <= 6'h00;
      write_address_data_log_force[8292] <= 6'h00;
      write_address_data_log_force[8293] <= 6'h00;
      write_address_data_log_force[8294] <= 6'h00;
      write_address_data_log_force[8295] <= 6'h00;
      write_address_data_log_force[8296] <= 6'h00;
      write_address_data_log_force[8297] <= 6'h00;
      write_address_data_log_force[8298] <= 6'h00;
      write_address_data_log_force[8299] <= 6'h00;
      write_address_data_log_force[8300] <= 6'h00;
      write_address_data_log_force[8301] <= 6'h00;
      write_address_data_log_force[8302] <= 6'h00;
      write_address_data_log_force[8303] <= 6'h00;
      write_address_data_log_force[8304] <= 6'h00;
      write_address_data_log_force[8305] <= 6'h00;
      write_address_data_log_force[8306] <= 6'h00;
      write_address_data_log_force[8307] <= 6'h00;
      write_address_data_log_force[8308] <= 6'h00;
      write_address_data_log_force[8309] <= 6'h00;
      write_address_data_log_force[8310] <= 6'h00;
      write_address_data_log_force[8311] <= 6'h00;
      write_address_data_log_force[8312] <= 6'h00;
      write_address_data_log_force[8313] <= 6'h00;
      write_address_data_log_force[8314] <= 6'h00;
      write_address_data_log_force[8315] <= 6'h00;
      write_address_data_log_force[8316] <= 6'h00;
      write_address_data_log_force[8317] <= 6'h00;
      write_address_data_log_force[8318] <= 6'h00;
      write_address_data_log_force[8319] <= 6'h00;

      // Input data for coeffs_in_data_log
      coeffs_in_data_log_force[   0] <= 16'hffd7;
      coeffs_in_data_log_force[   1] <= 16'hff83;
      coeffs_in_data_log_force[   2] <= 16'hff2e;
      coeffs_in_data_log_force[   3] <= 16'hfedf;
      coeffs_in_data_log_force[   4] <= 16'hfea6;
      coeffs_in_data_log_force[   5] <= 16'hfe9b;
      coeffs_in_data_log_force[   6] <= 16'hfedc;
      coeffs_in_data_log_force[   7] <= 16'hff83;
      coeffs_in_data_log_force[   8] <= 16'h0098;
      coeffs_in_data_log_force[   9] <= 16'h020b;
      coeffs_in_data_log_force[  10] <= 16'h03ac;
      coeffs_in_data_log_force[  11] <= 16'h0529;
      coeffs_in_data_log_force[  12] <= 16'h061d;
      coeffs_in_data_log_force[  13] <= 16'h061a;
      coeffs_in_data_log_force[  14] <= 16'h04c6;
      coeffs_in_data_log_force[  15] <= 16'h01f4;
      coeffs_in_data_log_force[  16] <= 16'hfdbb;
      coeffs_in_data_log_force[  17] <= 16'hf886;
      coeffs_in_data_log_force[  18] <= 16'hf312;
      coeffs_in_data_log_force[  19] <= 16'hee66;
      coeffs_in_data_log_force[  20] <= 16'hebad;
      coeffs_in_data_log_force[  21] <= 16'hec13;
      coeffs_in_data_log_force[  22] <= 16'hf08c;
      coeffs_in_data_log_force[  23] <= 16'hf9ab;
      coeffs_in_data_log_force[  24] <= 16'h0775;
      coeffs_in_data_log_force[  25] <= 16'h1953;
      coeffs_in_data_log_force[  26] <= 16'h2e12;
      coeffs_in_data_log_force[  27] <= 16'h43fc;
      coeffs_in_data_log_force[  28] <= 16'h590a;
      coeffs_in_data_log_force[  29] <= 16'h6b25;
      coeffs_in_data_log_force[  30] <= 16'h786c;
      coeffs_in_data_log_force[  31] <= 16'h7f71;
      coeffs_in_data_log_force[  32] <= 16'h7f71;
      coeffs_in_data_log_force[  33] <= 16'h786c;
      coeffs_in_data_log_force[  34] <= 16'h6b25;
      coeffs_in_data_log_force[  35] <= 16'h590a;
      coeffs_in_data_log_force[  36] <= 16'h43fc;
      coeffs_in_data_log_force[  37] <= 16'h2e12;
      coeffs_in_data_log_force[  38] <= 16'h1953;
      coeffs_in_data_log_force[  39] <= 16'h0775;
      coeffs_in_data_log_force[  40] <= 16'hf9ab;
      coeffs_in_data_log_force[  41] <= 16'hf08c;
      coeffs_in_data_log_force[  42] <= 16'hec13;
      coeffs_in_data_log_force[  43] <= 16'hebad;
      coeffs_in_data_log_force[  44] <= 16'hee66;
      coeffs_in_data_log_force[  45] <= 16'hf312;
      coeffs_in_data_log_force[  46] <= 16'hf886;
      coeffs_in_data_log_force[  47] <= 16'hfdbb;
      coeffs_in_data_log_force[  48] <= 16'h01f4;
      coeffs_in_data_log_force[  49] <= 16'h04c6;
      coeffs_in_data_log_force[  50] <= 16'h061a;
      coeffs_in_data_log_force[  51] <= 16'h061d;
      coeffs_in_data_log_force[  52] <= 16'h0529;
      coeffs_in_data_log_force[  53] <= 16'h03ac;
      coeffs_in_data_log_force[  54] <= 16'h020b;
      coeffs_in_data_log_force[  55] <= 16'h0098;
      coeffs_in_data_log_force[  56] <= 16'hff83;
      coeffs_in_data_log_force[  57] <= 16'hfedc;
      coeffs_in_data_log_force[  58] <= 16'hfe9b;
      coeffs_in_data_log_force[  59] <= 16'hfea6;
      coeffs_in_data_log_force[  60] <= 16'hfedf;
      coeffs_in_data_log_force[  61] <= 16'hff2e;
      coeffs_in_data_log_force[  62] <= 16'hff83;
      coeffs_in_data_log_force[  63] <= 16'hffd7;
      coeffs_in_data_log_force[  64] <= 16'h0000;
      coeffs_in_data_log_force[  65] <= 16'h0000;
      coeffs_in_data_log_force[  66] <= 16'h0000;
      coeffs_in_data_log_force[  67] <= 16'h0000;
      coeffs_in_data_log_force[  68] <= 16'h0000;
      coeffs_in_data_log_force[  69] <= 16'h0000;
      coeffs_in_data_log_force[  70] <= 16'h0000;
      coeffs_in_data_log_force[  71] <= 16'h0000;
      coeffs_in_data_log_force[  72] <= 16'h0000;
      coeffs_in_data_log_force[  73] <= 16'h0000;
      coeffs_in_data_log_force[  74] <= 16'h0000;
      coeffs_in_data_log_force[  75] <= 16'h0000;
      coeffs_in_data_log_force[  76] <= 16'h0000;
      coeffs_in_data_log_force[  77] <= 16'h0000;
      coeffs_in_data_log_force[  78] <= 16'h0000;
      coeffs_in_data_log_force[  79] <= 16'h0000;
      coeffs_in_data_log_force[  80] <= 16'h0000;
      coeffs_in_data_log_force[  81] <= 16'h0000;
      coeffs_in_data_log_force[  82] <= 16'h0000;
      coeffs_in_data_log_force[  83] <= 16'h0000;
      coeffs_in_data_log_force[  84] <= 16'h0000;
      coeffs_in_data_log_force[  85] <= 16'h0000;
      coeffs_in_data_log_force[  86] <= 16'h0000;
      coeffs_in_data_log_force[  87] <= 16'h0000;
      coeffs_in_data_log_force[  88] <= 16'h0000;
      coeffs_in_data_log_force[  89] <= 16'h0000;
      coeffs_in_data_log_force[  90] <= 16'h0000;
      coeffs_in_data_log_force[  91] <= 16'h0000;
      coeffs_in_data_log_force[  92] <= 16'h0000;
      coeffs_in_data_log_force[  93] <= 16'h0000;
      coeffs_in_data_log_force[  94] <= 16'h0000;
      coeffs_in_data_log_force[  95] <= 16'h0000;
      coeffs_in_data_log_force[  96] <= 16'h0000;
      coeffs_in_data_log_force[  97] <= 16'h0000;
      coeffs_in_data_log_force[  98] <= 16'h0000;
      coeffs_in_data_log_force[  99] <= 16'h0000;
      coeffs_in_data_log_force[ 100] <= 16'h0000;
      coeffs_in_data_log_force[ 101] <= 16'h0000;
      coeffs_in_data_log_force[ 102] <= 16'h0000;
      coeffs_in_data_log_force[ 103] <= 16'h0000;
      coeffs_in_data_log_force[ 104] <= 16'h0000;
      coeffs_in_data_log_force[ 105] <= 16'h0000;
      coeffs_in_data_log_force[ 106] <= 16'h0000;
      coeffs_in_data_log_force[ 107] <= 16'h0000;
      coeffs_in_data_log_force[ 108] <= 16'h0000;
      coeffs_in_data_log_force[ 109] <= 16'h0000;
      coeffs_in_data_log_force[ 110] <= 16'h0000;
      coeffs_in_data_log_force[ 111] <= 16'h0000;
      coeffs_in_data_log_force[ 112] <= 16'h0000;
      coeffs_in_data_log_force[ 113] <= 16'h0000;
      coeffs_in_data_log_force[ 114] <= 16'h0000;
      coeffs_in_data_log_force[ 115] <= 16'h0000;
      coeffs_in_data_log_force[ 116] <= 16'h0000;
      coeffs_in_data_log_force[ 117] <= 16'h0000;
      coeffs_in_data_log_force[ 118] <= 16'h0000;
      coeffs_in_data_log_force[ 119] <= 16'h0000;
      coeffs_in_data_log_force[ 120] <= 16'h0000;
      coeffs_in_data_log_force[ 121] <= 16'h0000;
      coeffs_in_data_log_force[ 122] <= 16'h0000;
      coeffs_in_data_log_force[ 123] <= 16'h0000;
      coeffs_in_data_log_force[ 124] <= 16'h0000;
      coeffs_in_data_log_force[ 125] <= 16'h0000;
      coeffs_in_data_log_force[ 126] <= 16'h0000;
      coeffs_in_data_log_force[ 127] <= 16'h0000;
      coeffs_in_data_log_force[ 128] <= 16'h0000;
      coeffs_in_data_log_force[ 129] <= 16'h0000;
      coeffs_in_data_log_force[ 130] <= 16'h0000;
      coeffs_in_data_log_force[ 131] <= 16'h0000;
      coeffs_in_data_log_force[ 132] <= 16'h0000;
      coeffs_in_data_log_force[ 133] <= 16'h0000;
      coeffs_in_data_log_force[ 134] <= 16'h0000;
      coeffs_in_data_log_force[ 135] <= 16'h0000;
      coeffs_in_data_log_force[ 136] <= 16'h0000;
      coeffs_in_data_log_force[ 137] <= 16'h0000;
      coeffs_in_data_log_force[ 138] <= 16'h0000;
      coeffs_in_data_log_force[ 139] <= 16'h0000;
      coeffs_in_data_log_force[ 140] <= 16'h0000;
      coeffs_in_data_log_force[ 141] <= 16'h0000;
      coeffs_in_data_log_force[ 142] <= 16'h0000;
      coeffs_in_data_log_force[ 143] <= 16'h0000;
      coeffs_in_data_log_force[ 144] <= 16'h0000;
      coeffs_in_data_log_force[ 145] <= 16'h0000;
      coeffs_in_data_log_force[ 146] <= 16'h0000;
      coeffs_in_data_log_force[ 147] <= 16'h0000;
      coeffs_in_data_log_force[ 148] <= 16'h0000;
      coeffs_in_data_log_force[ 149] <= 16'h0000;
      coeffs_in_data_log_force[ 150] <= 16'h0000;
      coeffs_in_data_log_force[ 151] <= 16'h0000;
      coeffs_in_data_log_force[ 152] <= 16'h0000;
      coeffs_in_data_log_force[ 153] <= 16'h0000;
      coeffs_in_data_log_force[ 154] <= 16'h0000;
      coeffs_in_data_log_force[ 155] <= 16'h0000;
      coeffs_in_data_log_force[ 156] <= 16'h0000;
      coeffs_in_data_log_force[ 157] <= 16'h0000;
      coeffs_in_data_log_force[ 158] <= 16'h0000;
      coeffs_in_data_log_force[ 159] <= 16'h0000;
      coeffs_in_data_log_force[ 160] <= 16'h0000;
      coeffs_in_data_log_force[ 161] <= 16'h0000;
      coeffs_in_data_log_force[ 162] <= 16'h0000;
      coeffs_in_data_log_force[ 163] <= 16'h0000;
      coeffs_in_data_log_force[ 164] <= 16'h0000;
      coeffs_in_data_log_force[ 165] <= 16'h0000;
      coeffs_in_data_log_force[ 166] <= 16'h0000;
      coeffs_in_data_log_force[ 167] <= 16'h0000;
      coeffs_in_data_log_force[ 168] <= 16'h0000;
      coeffs_in_data_log_force[ 169] <= 16'h0000;
      coeffs_in_data_log_force[ 170] <= 16'h0000;
      coeffs_in_data_log_force[ 171] <= 16'h0000;
      coeffs_in_data_log_force[ 172] <= 16'h0000;
      coeffs_in_data_log_force[ 173] <= 16'h0000;
      coeffs_in_data_log_force[ 174] <= 16'h0000;
      coeffs_in_data_log_force[ 175] <= 16'h0000;
      coeffs_in_data_log_force[ 176] <= 16'h0000;
      coeffs_in_data_log_force[ 177] <= 16'h0000;
      coeffs_in_data_log_force[ 178] <= 16'h0000;
      coeffs_in_data_log_force[ 179] <= 16'h0000;
      coeffs_in_data_log_force[ 180] <= 16'h0000;
      coeffs_in_data_log_force[ 181] <= 16'h0000;
      coeffs_in_data_log_force[ 182] <= 16'h0000;
      coeffs_in_data_log_force[ 183] <= 16'h0000;
      coeffs_in_data_log_force[ 184] <= 16'h0000;
      coeffs_in_data_log_force[ 185] <= 16'h0000;
      coeffs_in_data_log_force[ 186] <= 16'h0000;
      coeffs_in_data_log_force[ 187] <= 16'h0000;
      coeffs_in_data_log_force[ 188] <= 16'h0000;
      coeffs_in_data_log_force[ 189] <= 16'h0000;
      coeffs_in_data_log_force[ 190] <= 16'h0000;
      coeffs_in_data_log_force[ 191] <= 16'h0000;
      coeffs_in_data_log_force[ 192] <= 16'h0000;
      coeffs_in_data_log_force[ 193] <= 16'h0000;
      coeffs_in_data_log_force[ 194] <= 16'h0000;
      coeffs_in_data_log_force[ 195] <= 16'h0000;
      coeffs_in_data_log_force[ 196] <= 16'h0000;
      coeffs_in_data_log_force[ 197] <= 16'h0000;
      coeffs_in_data_log_force[ 198] <= 16'h0000;
      coeffs_in_data_log_force[ 199] <= 16'h0000;
      coeffs_in_data_log_force[ 200] <= 16'h0000;
      coeffs_in_data_log_force[ 201] <= 16'h0000;
      coeffs_in_data_log_force[ 202] <= 16'h0000;
      coeffs_in_data_log_force[ 203] <= 16'h0000;
      coeffs_in_data_log_force[ 204] <= 16'h0000;
      coeffs_in_data_log_force[ 205] <= 16'h0000;
      coeffs_in_data_log_force[ 206] <= 16'h0000;
      coeffs_in_data_log_force[ 207] <= 16'h0000;
      coeffs_in_data_log_force[ 208] <= 16'h0000;
      coeffs_in_data_log_force[ 209] <= 16'h0000;
      coeffs_in_data_log_force[ 210] <= 16'h0000;
      coeffs_in_data_log_force[ 211] <= 16'h0000;
      coeffs_in_data_log_force[ 212] <= 16'h0000;
      coeffs_in_data_log_force[ 213] <= 16'h0000;
      coeffs_in_data_log_force[ 214] <= 16'h0000;
      coeffs_in_data_log_force[ 215] <= 16'h0000;
      coeffs_in_data_log_force[ 216] <= 16'h0000;
      coeffs_in_data_log_force[ 217] <= 16'h0000;
      coeffs_in_data_log_force[ 218] <= 16'h0000;
      coeffs_in_data_log_force[ 219] <= 16'h0000;
      coeffs_in_data_log_force[ 220] <= 16'h0000;
      coeffs_in_data_log_force[ 221] <= 16'h0000;
      coeffs_in_data_log_force[ 222] <= 16'h0000;
      coeffs_in_data_log_force[ 223] <= 16'h0000;
      coeffs_in_data_log_force[ 224] <= 16'h0000;
      coeffs_in_data_log_force[ 225] <= 16'h0000;
      coeffs_in_data_log_force[ 226] <= 16'h0000;
      coeffs_in_data_log_force[ 227] <= 16'h0000;
      coeffs_in_data_log_force[ 228] <= 16'h0000;
      coeffs_in_data_log_force[ 229] <= 16'h0000;
      coeffs_in_data_log_force[ 230] <= 16'h0000;
      coeffs_in_data_log_force[ 231] <= 16'h0000;
      coeffs_in_data_log_force[ 232] <= 16'h0000;
      coeffs_in_data_log_force[ 233] <= 16'h0000;
      coeffs_in_data_log_force[ 234] <= 16'h0000;
      coeffs_in_data_log_force[ 235] <= 16'h0000;
      coeffs_in_data_log_force[ 236] <= 16'h0000;
      coeffs_in_data_log_force[ 237] <= 16'h0000;
      coeffs_in_data_log_force[ 238] <= 16'h0000;
      coeffs_in_data_log_force[ 239] <= 16'h0000;
      coeffs_in_data_log_force[ 240] <= 16'h0000;
      coeffs_in_data_log_force[ 241] <= 16'h0000;
      coeffs_in_data_log_force[ 242] <= 16'h0000;
      coeffs_in_data_log_force[ 243] <= 16'h0000;
      coeffs_in_data_log_force[ 244] <= 16'h0000;
      coeffs_in_data_log_force[ 245] <= 16'h0000;
      coeffs_in_data_log_force[ 246] <= 16'h0000;
      coeffs_in_data_log_force[ 247] <= 16'h0000;
      coeffs_in_data_log_force[ 248] <= 16'h0000;
      coeffs_in_data_log_force[ 249] <= 16'h0000;
      coeffs_in_data_log_force[ 250] <= 16'h0000;
      coeffs_in_data_log_force[ 251] <= 16'h0000;
      coeffs_in_data_log_force[ 252] <= 16'h0000;
      coeffs_in_data_log_force[ 253] <= 16'h0000;
      coeffs_in_data_log_force[ 254] <= 16'h0000;
      coeffs_in_data_log_force[ 255] <= 16'h0000;
      coeffs_in_data_log_force[ 256] <= 16'h0000;
      coeffs_in_data_log_force[ 257] <= 16'h0000;
      coeffs_in_data_log_force[ 258] <= 16'h0000;
      coeffs_in_data_log_force[ 259] <= 16'h0000;
      coeffs_in_data_log_force[ 260] <= 16'h0000;
      coeffs_in_data_log_force[ 261] <= 16'h0000;
      coeffs_in_data_log_force[ 262] <= 16'h0000;
      coeffs_in_data_log_force[ 263] <= 16'h0000;
      coeffs_in_data_log_force[ 264] <= 16'h0000;
      coeffs_in_data_log_force[ 265] <= 16'h0000;
      coeffs_in_data_log_force[ 266] <= 16'h0000;
      coeffs_in_data_log_force[ 267] <= 16'h0000;
      coeffs_in_data_log_force[ 268] <= 16'h0000;
      coeffs_in_data_log_force[ 269] <= 16'h0000;
      coeffs_in_data_log_force[ 270] <= 16'h0000;
      coeffs_in_data_log_force[ 271] <= 16'h0000;
      coeffs_in_data_log_force[ 272] <= 16'h0000;
      coeffs_in_data_log_force[ 273] <= 16'h0000;
      coeffs_in_data_log_force[ 274] <= 16'h0000;
      coeffs_in_data_log_force[ 275] <= 16'h0000;
      coeffs_in_data_log_force[ 276] <= 16'h0000;
      coeffs_in_data_log_force[ 277] <= 16'h0000;
      coeffs_in_data_log_force[ 278] <= 16'h0000;
      coeffs_in_data_log_force[ 279] <= 16'h0000;
      coeffs_in_data_log_force[ 280] <= 16'h0000;
      coeffs_in_data_log_force[ 281] <= 16'h0000;
      coeffs_in_data_log_force[ 282] <= 16'h0000;
      coeffs_in_data_log_force[ 283] <= 16'h0000;
      coeffs_in_data_log_force[ 284] <= 16'h0000;
      coeffs_in_data_log_force[ 285] <= 16'h0000;
      coeffs_in_data_log_force[ 286] <= 16'h0000;
      coeffs_in_data_log_force[ 287] <= 16'h0000;
      coeffs_in_data_log_force[ 288] <= 16'h0000;
      coeffs_in_data_log_force[ 289] <= 16'h0000;
      coeffs_in_data_log_force[ 290] <= 16'h0000;
      coeffs_in_data_log_force[ 291] <= 16'h0000;
      coeffs_in_data_log_force[ 292] <= 16'h0000;
      coeffs_in_data_log_force[ 293] <= 16'h0000;
      coeffs_in_data_log_force[ 294] <= 16'h0000;
      coeffs_in_data_log_force[ 295] <= 16'h0000;
      coeffs_in_data_log_force[ 296] <= 16'h0000;
      coeffs_in_data_log_force[ 297] <= 16'h0000;
      coeffs_in_data_log_force[ 298] <= 16'h0000;
      coeffs_in_data_log_force[ 299] <= 16'h0000;
      coeffs_in_data_log_force[ 300] <= 16'h0000;
      coeffs_in_data_log_force[ 301] <= 16'h0000;
      coeffs_in_data_log_force[ 302] <= 16'h0000;
      coeffs_in_data_log_force[ 303] <= 16'h0000;
      coeffs_in_data_log_force[ 304] <= 16'h0000;
      coeffs_in_data_log_force[ 305] <= 16'h0000;
      coeffs_in_data_log_force[ 306] <= 16'h0000;
      coeffs_in_data_log_force[ 307] <= 16'h0000;
      coeffs_in_data_log_force[ 308] <= 16'h0000;
      coeffs_in_data_log_force[ 309] <= 16'h0000;
      coeffs_in_data_log_force[ 310] <= 16'h0000;
      coeffs_in_data_log_force[ 311] <= 16'h0000;
      coeffs_in_data_log_force[ 312] <= 16'h0000;
      coeffs_in_data_log_force[ 313] <= 16'h0000;
      coeffs_in_data_log_force[ 314] <= 16'h0000;
      coeffs_in_data_log_force[ 315] <= 16'h0000;
      coeffs_in_data_log_force[ 316] <= 16'h0000;
      coeffs_in_data_log_force[ 317] <= 16'h0000;
      coeffs_in_data_log_force[ 318] <= 16'h0000;
      coeffs_in_data_log_force[ 319] <= 16'h0000;
      coeffs_in_data_log_force[ 320] <= 16'h0000;
      coeffs_in_data_log_force[ 321] <= 16'h0000;
      coeffs_in_data_log_force[ 322] <= 16'h0000;
      coeffs_in_data_log_force[ 323] <= 16'h0000;
      coeffs_in_data_log_force[ 324] <= 16'h0000;
      coeffs_in_data_log_force[ 325] <= 16'h0000;
      coeffs_in_data_log_force[ 326] <= 16'h0000;
      coeffs_in_data_log_force[ 327] <= 16'h0000;
      coeffs_in_data_log_force[ 328] <= 16'h0000;
      coeffs_in_data_log_force[ 329] <= 16'h0000;
      coeffs_in_data_log_force[ 330] <= 16'h0000;
      coeffs_in_data_log_force[ 331] <= 16'h0000;
      coeffs_in_data_log_force[ 332] <= 16'h0000;
      coeffs_in_data_log_force[ 333] <= 16'h0000;
      coeffs_in_data_log_force[ 334] <= 16'h0000;
      coeffs_in_data_log_force[ 335] <= 16'h0000;
      coeffs_in_data_log_force[ 336] <= 16'h0000;
      coeffs_in_data_log_force[ 337] <= 16'h0000;
      coeffs_in_data_log_force[ 338] <= 16'h0000;
      coeffs_in_data_log_force[ 339] <= 16'h0000;
      coeffs_in_data_log_force[ 340] <= 16'h0000;
      coeffs_in_data_log_force[ 341] <= 16'h0000;
      coeffs_in_data_log_force[ 342] <= 16'h0000;
      coeffs_in_data_log_force[ 343] <= 16'h0000;
      coeffs_in_data_log_force[ 344] <= 16'h0000;
      coeffs_in_data_log_force[ 345] <= 16'h0000;
      coeffs_in_data_log_force[ 346] <= 16'h0000;
      coeffs_in_data_log_force[ 347] <= 16'h0000;
      coeffs_in_data_log_force[ 348] <= 16'h0000;
      coeffs_in_data_log_force[ 349] <= 16'h0000;
      coeffs_in_data_log_force[ 350] <= 16'h0000;
      coeffs_in_data_log_force[ 351] <= 16'h0000;
      coeffs_in_data_log_force[ 352] <= 16'h0000;
      coeffs_in_data_log_force[ 353] <= 16'h0000;
      coeffs_in_data_log_force[ 354] <= 16'h0000;
      coeffs_in_data_log_force[ 355] <= 16'h0000;
      coeffs_in_data_log_force[ 356] <= 16'h0000;
      coeffs_in_data_log_force[ 357] <= 16'h0000;
      coeffs_in_data_log_force[ 358] <= 16'h0000;
      coeffs_in_data_log_force[ 359] <= 16'h0000;
      coeffs_in_data_log_force[ 360] <= 16'h0000;
      coeffs_in_data_log_force[ 361] <= 16'h0000;
      coeffs_in_data_log_force[ 362] <= 16'h0000;
      coeffs_in_data_log_force[ 363] <= 16'h0000;
      coeffs_in_data_log_force[ 364] <= 16'h0000;
      coeffs_in_data_log_force[ 365] <= 16'h0000;
      coeffs_in_data_log_force[ 366] <= 16'h0000;
      coeffs_in_data_log_force[ 367] <= 16'h0000;
      coeffs_in_data_log_force[ 368] <= 16'h0000;
      coeffs_in_data_log_force[ 369] <= 16'h0000;
      coeffs_in_data_log_force[ 370] <= 16'h0000;
      coeffs_in_data_log_force[ 371] <= 16'h0000;
      coeffs_in_data_log_force[ 372] <= 16'h0000;
      coeffs_in_data_log_force[ 373] <= 16'h0000;
      coeffs_in_data_log_force[ 374] <= 16'h0000;
      coeffs_in_data_log_force[ 375] <= 16'h0000;
      coeffs_in_data_log_force[ 376] <= 16'h0000;
      coeffs_in_data_log_force[ 377] <= 16'h0000;
      coeffs_in_data_log_force[ 378] <= 16'h0000;
      coeffs_in_data_log_force[ 379] <= 16'h0000;
      coeffs_in_data_log_force[ 380] <= 16'h0000;
      coeffs_in_data_log_force[ 381] <= 16'h0000;
      coeffs_in_data_log_force[ 382] <= 16'h0000;
      coeffs_in_data_log_force[ 383] <= 16'h0000;
      coeffs_in_data_log_force[ 384] <= 16'h0000;
      coeffs_in_data_log_force[ 385] <= 16'h0000;
      coeffs_in_data_log_force[ 386] <= 16'h0000;
      coeffs_in_data_log_force[ 387] <= 16'h0000;
      coeffs_in_data_log_force[ 388] <= 16'h0000;
      coeffs_in_data_log_force[ 389] <= 16'h0000;
      coeffs_in_data_log_force[ 390] <= 16'h0000;
      coeffs_in_data_log_force[ 391] <= 16'h0000;
      coeffs_in_data_log_force[ 392] <= 16'h0000;
      coeffs_in_data_log_force[ 393] <= 16'h0000;
      coeffs_in_data_log_force[ 394] <= 16'h0000;
      coeffs_in_data_log_force[ 395] <= 16'h0000;
      coeffs_in_data_log_force[ 396] <= 16'h0000;
      coeffs_in_data_log_force[ 397] <= 16'h0000;
      coeffs_in_data_log_force[ 398] <= 16'h0000;
      coeffs_in_data_log_force[ 399] <= 16'h0000;
      coeffs_in_data_log_force[ 400] <= 16'h0000;
      coeffs_in_data_log_force[ 401] <= 16'h0000;
      coeffs_in_data_log_force[ 402] <= 16'h0000;
      coeffs_in_data_log_force[ 403] <= 16'h0000;
      coeffs_in_data_log_force[ 404] <= 16'h0000;
      coeffs_in_data_log_force[ 405] <= 16'h0000;
      coeffs_in_data_log_force[ 406] <= 16'h0000;
      coeffs_in_data_log_force[ 407] <= 16'h0000;
      coeffs_in_data_log_force[ 408] <= 16'h0000;
      coeffs_in_data_log_force[ 409] <= 16'h0000;
      coeffs_in_data_log_force[ 410] <= 16'h0000;
      coeffs_in_data_log_force[ 411] <= 16'h0000;
      coeffs_in_data_log_force[ 412] <= 16'h0000;
      coeffs_in_data_log_force[ 413] <= 16'h0000;
      coeffs_in_data_log_force[ 414] <= 16'h0000;
      coeffs_in_data_log_force[ 415] <= 16'h0000;
      coeffs_in_data_log_force[ 416] <= 16'h0000;
      coeffs_in_data_log_force[ 417] <= 16'h0000;
      coeffs_in_data_log_force[ 418] <= 16'h0000;
      coeffs_in_data_log_force[ 419] <= 16'h0000;
      coeffs_in_data_log_force[ 420] <= 16'h0000;
      coeffs_in_data_log_force[ 421] <= 16'h0000;
      coeffs_in_data_log_force[ 422] <= 16'h0000;
      coeffs_in_data_log_force[ 423] <= 16'h0000;
      coeffs_in_data_log_force[ 424] <= 16'h0000;
      coeffs_in_data_log_force[ 425] <= 16'h0000;
      coeffs_in_data_log_force[ 426] <= 16'h0000;
      coeffs_in_data_log_force[ 427] <= 16'h0000;
      coeffs_in_data_log_force[ 428] <= 16'h0000;
      coeffs_in_data_log_force[ 429] <= 16'h0000;
      coeffs_in_data_log_force[ 430] <= 16'h0000;
      coeffs_in_data_log_force[ 431] <= 16'h0000;
      coeffs_in_data_log_force[ 432] <= 16'h0000;
      coeffs_in_data_log_force[ 433] <= 16'h0000;
      coeffs_in_data_log_force[ 434] <= 16'h0000;
      coeffs_in_data_log_force[ 435] <= 16'h0000;
      coeffs_in_data_log_force[ 436] <= 16'h0000;
      coeffs_in_data_log_force[ 437] <= 16'h0000;
      coeffs_in_data_log_force[ 438] <= 16'h0000;
      coeffs_in_data_log_force[ 439] <= 16'h0000;
      coeffs_in_data_log_force[ 440] <= 16'h0000;
      coeffs_in_data_log_force[ 441] <= 16'h0000;
      coeffs_in_data_log_force[ 442] <= 16'h0000;
      coeffs_in_data_log_force[ 443] <= 16'h0000;
      coeffs_in_data_log_force[ 444] <= 16'h0000;
      coeffs_in_data_log_force[ 445] <= 16'h0000;
      coeffs_in_data_log_force[ 446] <= 16'h0000;
      coeffs_in_data_log_force[ 447] <= 16'h0000;
      coeffs_in_data_log_force[ 448] <= 16'h0000;
      coeffs_in_data_log_force[ 449] <= 16'h0000;
      coeffs_in_data_log_force[ 450] <= 16'h0000;
      coeffs_in_data_log_force[ 451] <= 16'h0000;
      coeffs_in_data_log_force[ 452] <= 16'h0000;
      coeffs_in_data_log_force[ 453] <= 16'h0000;
      coeffs_in_data_log_force[ 454] <= 16'h0000;
      coeffs_in_data_log_force[ 455] <= 16'h0000;
      coeffs_in_data_log_force[ 456] <= 16'h0000;
      coeffs_in_data_log_force[ 457] <= 16'h0000;
      coeffs_in_data_log_force[ 458] <= 16'h0000;
      coeffs_in_data_log_force[ 459] <= 16'h0000;
      coeffs_in_data_log_force[ 460] <= 16'h0000;
      coeffs_in_data_log_force[ 461] <= 16'h0000;
      coeffs_in_data_log_force[ 462] <= 16'h0000;
      coeffs_in_data_log_force[ 463] <= 16'h0000;
      coeffs_in_data_log_force[ 464] <= 16'h0000;
      coeffs_in_data_log_force[ 465] <= 16'h0000;
      coeffs_in_data_log_force[ 466] <= 16'h0000;
      coeffs_in_data_log_force[ 467] <= 16'h0000;
      coeffs_in_data_log_force[ 468] <= 16'h0000;
      coeffs_in_data_log_force[ 469] <= 16'h0000;
      coeffs_in_data_log_force[ 470] <= 16'h0000;
      coeffs_in_data_log_force[ 471] <= 16'h0000;
      coeffs_in_data_log_force[ 472] <= 16'h0000;
      coeffs_in_data_log_force[ 473] <= 16'h0000;
      coeffs_in_data_log_force[ 474] <= 16'h0000;
      coeffs_in_data_log_force[ 475] <= 16'h0000;
      coeffs_in_data_log_force[ 476] <= 16'h0000;
      coeffs_in_data_log_force[ 477] <= 16'h0000;
      coeffs_in_data_log_force[ 478] <= 16'h0000;
      coeffs_in_data_log_force[ 479] <= 16'h0000;
      coeffs_in_data_log_force[ 480] <= 16'h0000;
      coeffs_in_data_log_force[ 481] <= 16'h0000;
      coeffs_in_data_log_force[ 482] <= 16'h0000;
      coeffs_in_data_log_force[ 483] <= 16'h0000;
      coeffs_in_data_log_force[ 484] <= 16'h0000;
      coeffs_in_data_log_force[ 485] <= 16'h0000;
      coeffs_in_data_log_force[ 486] <= 16'h0000;
      coeffs_in_data_log_force[ 487] <= 16'h0000;
      coeffs_in_data_log_force[ 488] <= 16'h0000;
      coeffs_in_data_log_force[ 489] <= 16'h0000;
      coeffs_in_data_log_force[ 490] <= 16'h0000;
      coeffs_in_data_log_force[ 491] <= 16'h0000;
      coeffs_in_data_log_force[ 492] <= 16'h0000;
      coeffs_in_data_log_force[ 493] <= 16'h0000;
      coeffs_in_data_log_force[ 494] <= 16'h0000;
      coeffs_in_data_log_force[ 495] <= 16'h0000;
      coeffs_in_data_log_force[ 496] <= 16'h0000;
      coeffs_in_data_log_force[ 497] <= 16'h0000;
      coeffs_in_data_log_force[ 498] <= 16'h0000;
      coeffs_in_data_log_force[ 499] <= 16'h0000;
      coeffs_in_data_log_force[ 500] <= 16'h0000;
      coeffs_in_data_log_force[ 501] <= 16'h0000;
      coeffs_in_data_log_force[ 502] <= 16'h0000;
      coeffs_in_data_log_force[ 503] <= 16'h0000;
      coeffs_in_data_log_force[ 504] <= 16'h0000;
      coeffs_in_data_log_force[ 505] <= 16'h0000;
      coeffs_in_data_log_force[ 506] <= 16'h0000;
      coeffs_in_data_log_force[ 507] <= 16'h0000;
      coeffs_in_data_log_force[ 508] <= 16'h0000;
      coeffs_in_data_log_force[ 509] <= 16'h0000;
      coeffs_in_data_log_force[ 510] <= 16'h0000;
      coeffs_in_data_log_force[ 511] <= 16'h0000;
      coeffs_in_data_log_force[ 512] <= 16'h0000;
      coeffs_in_data_log_force[ 513] <= 16'h0000;
      coeffs_in_data_log_force[ 514] <= 16'h0000;
      coeffs_in_data_log_force[ 515] <= 16'h0000;
      coeffs_in_data_log_force[ 516] <= 16'h0000;
      coeffs_in_data_log_force[ 517] <= 16'h0000;
      coeffs_in_data_log_force[ 518] <= 16'h0000;
      coeffs_in_data_log_force[ 519] <= 16'h0000;
      coeffs_in_data_log_force[ 520] <= 16'h0000;
      coeffs_in_data_log_force[ 521] <= 16'h0000;
      coeffs_in_data_log_force[ 522] <= 16'h0000;
      coeffs_in_data_log_force[ 523] <= 16'h0000;
      coeffs_in_data_log_force[ 524] <= 16'h0000;
      coeffs_in_data_log_force[ 525] <= 16'h0000;
      coeffs_in_data_log_force[ 526] <= 16'h0000;
      coeffs_in_data_log_force[ 527] <= 16'h0000;
      coeffs_in_data_log_force[ 528] <= 16'h0000;
      coeffs_in_data_log_force[ 529] <= 16'h0000;
      coeffs_in_data_log_force[ 530] <= 16'h0000;
      coeffs_in_data_log_force[ 531] <= 16'h0000;
      coeffs_in_data_log_force[ 532] <= 16'h0000;
      coeffs_in_data_log_force[ 533] <= 16'h0000;
      coeffs_in_data_log_force[ 534] <= 16'h0000;
      coeffs_in_data_log_force[ 535] <= 16'h0000;
      coeffs_in_data_log_force[ 536] <= 16'h0000;
      coeffs_in_data_log_force[ 537] <= 16'h0000;
      coeffs_in_data_log_force[ 538] <= 16'h0000;
      coeffs_in_data_log_force[ 539] <= 16'h0000;
      coeffs_in_data_log_force[ 540] <= 16'h0000;
      coeffs_in_data_log_force[ 541] <= 16'h0000;
      coeffs_in_data_log_force[ 542] <= 16'h0000;
      coeffs_in_data_log_force[ 543] <= 16'h0000;
      coeffs_in_data_log_force[ 544] <= 16'h0000;
      coeffs_in_data_log_force[ 545] <= 16'h0000;
      coeffs_in_data_log_force[ 546] <= 16'h0000;
      coeffs_in_data_log_force[ 547] <= 16'h0000;
      coeffs_in_data_log_force[ 548] <= 16'h0000;
      coeffs_in_data_log_force[ 549] <= 16'h0000;
      coeffs_in_data_log_force[ 550] <= 16'h0000;
      coeffs_in_data_log_force[ 551] <= 16'h0000;
      coeffs_in_data_log_force[ 552] <= 16'h0000;
      coeffs_in_data_log_force[ 553] <= 16'h0000;
      coeffs_in_data_log_force[ 554] <= 16'h0000;
      coeffs_in_data_log_force[ 555] <= 16'h0000;
      coeffs_in_data_log_force[ 556] <= 16'h0000;
      coeffs_in_data_log_force[ 557] <= 16'h0000;
      coeffs_in_data_log_force[ 558] <= 16'h0000;
      coeffs_in_data_log_force[ 559] <= 16'h0000;
      coeffs_in_data_log_force[ 560] <= 16'h0000;
      coeffs_in_data_log_force[ 561] <= 16'h0000;
      coeffs_in_data_log_force[ 562] <= 16'h0000;
      coeffs_in_data_log_force[ 563] <= 16'h0000;
      coeffs_in_data_log_force[ 564] <= 16'h0000;
      coeffs_in_data_log_force[ 565] <= 16'h0000;
      coeffs_in_data_log_force[ 566] <= 16'h0000;
      coeffs_in_data_log_force[ 567] <= 16'h0000;
      coeffs_in_data_log_force[ 568] <= 16'h0000;
      coeffs_in_data_log_force[ 569] <= 16'h0000;
      coeffs_in_data_log_force[ 570] <= 16'h0000;
      coeffs_in_data_log_force[ 571] <= 16'h0000;
      coeffs_in_data_log_force[ 572] <= 16'h0000;
      coeffs_in_data_log_force[ 573] <= 16'h0000;
      coeffs_in_data_log_force[ 574] <= 16'h0000;
      coeffs_in_data_log_force[ 575] <= 16'h0000;
      coeffs_in_data_log_force[ 576] <= 16'h0000;
      coeffs_in_data_log_force[ 577] <= 16'h0000;
      coeffs_in_data_log_force[ 578] <= 16'h0000;
      coeffs_in_data_log_force[ 579] <= 16'h0000;
      coeffs_in_data_log_force[ 580] <= 16'h0000;
      coeffs_in_data_log_force[ 581] <= 16'h0000;
      coeffs_in_data_log_force[ 582] <= 16'h0000;
      coeffs_in_data_log_force[ 583] <= 16'h0000;
      coeffs_in_data_log_force[ 584] <= 16'h0000;
      coeffs_in_data_log_force[ 585] <= 16'h0000;
      coeffs_in_data_log_force[ 586] <= 16'h0000;
      coeffs_in_data_log_force[ 587] <= 16'h0000;
      coeffs_in_data_log_force[ 588] <= 16'h0000;
      coeffs_in_data_log_force[ 589] <= 16'h0000;
      coeffs_in_data_log_force[ 590] <= 16'h0000;
      coeffs_in_data_log_force[ 591] <= 16'h0000;
      coeffs_in_data_log_force[ 592] <= 16'h0000;
      coeffs_in_data_log_force[ 593] <= 16'h0000;
      coeffs_in_data_log_force[ 594] <= 16'h0000;
      coeffs_in_data_log_force[ 595] <= 16'h0000;
      coeffs_in_data_log_force[ 596] <= 16'h0000;
      coeffs_in_data_log_force[ 597] <= 16'h0000;
      coeffs_in_data_log_force[ 598] <= 16'h0000;
      coeffs_in_data_log_force[ 599] <= 16'h0000;
      coeffs_in_data_log_force[ 600] <= 16'h0000;
      coeffs_in_data_log_force[ 601] <= 16'h0000;
      coeffs_in_data_log_force[ 602] <= 16'h0000;
      coeffs_in_data_log_force[ 603] <= 16'h0000;
      coeffs_in_data_log_force[ 604] <= 16'h0000;
      coeffs_in_data_log_force[ 605] <= 16'h0000;
      coeffs_in_data_log_force[ 606] <= 16'h0000;
      coeffs_in_data_log_force[ 607] <= 16'h0000;
      coeffs_in_data_log_force[ 608] <= 16'h0000;
      coeffs_in_data_log_force[ 609] <= 16'h0000;
      coeffs_in_data_log_force[ 610] <= 16'h0000;
      coeffs_in_data_log_force[ 611] <= 16'h0000;
      coeffs_in_data_log_force[ 612] <= 16'h0000;
      coeffs_in_data_log_force[ 613] <= 16'h0000;
      coeffs_in_data_log_force[ 614] <= 16'h0000;
      coeffs_in_data_log_force[ 615] <= 16'h0000;
      coeffs_in_data_log_force[ 616] <= 16'h0000;
      coeffs_in_data_log_force[ 617] <= 16'h0000;
      coeffs_in_data_log_force[ 618] <= 16'h0000;
      coeffs_in_data_log_force[ 619] <= 16'h0000;
      coeffs_in_data_log_force[ 620] <= 16'h0000;
      coeffs_in_data_log_force[ 621] <= 16'h0000;
      coeffs_in_data_log_force[ 622] <= 16'h0000;
      coeffs_in_data_log_force[ 623] <= 16'h0000;
      coeffs_in_data_log_force[ 624] <= 16'h0000;
      coeffs_in_data_log_force[ 625] <= 16'h0000;
      coeffs_in_data_log_force[ 626] <= 16'h0000;
      coeffs_in_data_log_force[ 627] <= 16'h0000;
      coeffs_in_data_log_force[ 628] <= 16'h0000;
      coeffs_in_data_log_force[ 629] <= 16'h0000;
      coeffs_in_data_log_force[ 630] <= 16'h0000;
      coeffs_in_data_log_force[ 631] <= 16'h0000;
      coeffs_in_data_log_force[ 632] <= 16'h0000;
      coeffs_in_data_log_force[ 633] <= 16'h0000;
      coeffs_in_data_log_force[ 634] <= 16'h0000;
      coeffs_in_data_log_force[ 635] <= 16'h0000;
      coeffs_in_data_log_force[ 636] <= 16'h0000;
      coeffs_in_data_log_force[ 637] <= 16'h0000;
      coeffs_in_data_log_force[ 638] <= 16'h0000;
      coeffs_in_data_log_force[ 639] <= 16'h0000;
      coeffs_in_data_log_force[ 640] <= 16'h0000;
      coeffs_in_data_log_force[ 641] <= 16'h0000;
      coeffs_in_data_log_force[ 642] <= 16'h0000;
      coeffs_in_data_log_force[ 643] <= 16'h0000;
      coeffs_in_data_log_force[ 644] <= 16'h0000;
      coeffs_in_data_log_force[ 645] <= 16'h0000;
      coeffs_in_data_log_force[ 646] <= 16'h0000;
      coeffs_in_data_log_force[ 647] <= 16'h0000;
      coeffs_in_data_log_force[ 648] <= 16'h0000;
      coeffs_in_data_log_force[ 649] <= 16'h0000;
      coeffs_in_data_log_force[ 650] <= 16'h0000;
      coeffs_in_data_log_force[ 651] <= 16'h0000;
      coeffs_in_data_log_force[ 652] <= 16'h0000;
      coeffs_in_data_log_force[ 653] <= 16'h0000;
      coeffs_in_data_log_force[ 654] <= 16'h0000;
      coeffs_in_data_log_force[ 655] <= 16'h0000;
      coeffs_in_data_log_force[ 656] <= 16'h0000;
      coeffs_in_data_log_force[ 657] <= 16'h0000;
      coeffs_in_data_log_force[ 658] <= 16'h0000;
      coeffs_in_data_log_force[ 659] <= 16'h0000;
      coeffs_in_data_log_force[ 660] <= 16'h0000;
      coeffs_in_data_log_force[ 661] <= 16'h0000;
      coeffs_in_data_log_force[ 662] <= 16'h0000;
      coeffs_in_data_log_force[ 663] <= 16'h0000;
      coeffs_in_data_log_force[ 664] <= 16'h0000;
      coeffs_in_data_log_force[ 665] <= 16'h0000;
      coeffs_in_data_log_force[ 666] <= 16'h0000;
      coeffs_in_data_log_force[ 667] <= 16'h0000;
      coeffs_in_data_log_force[ 668] <= 16'h0000;
      coeffs_in_data_log_force[ 669] <= 16'h0000;
      coeffs_in_data_log_force[ 670] <= 16'h0000;
      coeffs_in_data_log_force[ 671] <= 16'h0000;
      coeffs_in_data_log_force[ 672] <= 16'h0000;
      coeffs_in_data_log_force[ 673] <= 16'h0000;
      coeffs_in_data_log_force[ 674] <= 16'h0000;
      coeffs_in_data_log_force[ 675] <= 16'h0000;
      coeffs_in_data_log_force[ 676] <= 16'h0000;
      coeffs_in_data_log_force[ 677] <= 16'h0000;
      coeffs_in_data_log_force[ 678] <= 16'h0000;
      coeffs_in_data_log_force[ 679] <= 16'h0000;
      coeffs_in_data_log_force[ 680] <= 16'h0000;
      coeffs_in_data_log_force[ 681] <= 16'h0000;
      coeffs_in_data_log_force[ 682] <= 16'h0000;
      coeffs_in_data_log_force[ 683] <= 16'h0000;
      coeffs_in_data_log_force[ 684] <= 16'h0000;
      coeffs_in_data_log_force[ 685] <= 16'h0000;
      coeffs_in_data_log_force[ 686] <= 16'h0000;
      coeffs_in_data_log_force[ 687] <= 16'h0000;
      coeffs_in_data_log_force[ 688] <= 16'h0000;
      coeffs_in_data_log_force[ 689] <= 16'h0000;
      coeffs_in_data_log_force[ 690] <= 16'h0000;
      coeffs_in_data_log_force[ 691] <= 16'h0000;
      coeffs_in_data_log_force[ 692] <= 16'h0000;
      coeffs_in_data_log_force[ 693] <= 16'h0000;
      coeffs_in_data_log_force[ 694] <= 16'h0000;
      coeffs_in_data_log_force[ 695] <= 16'h0000;
      coeffs_in_data_log_force[ 696] <= 16'h0000;
      coeffs_in_data_log_force[ 697] <= 16'h0000;
      coeffs_in_data_log_force[ 698] <= 16'h0000;
      coeffs_in_data_log_force[ 699] <= 16'h0000;
      coeffs_in_data_log_force[ 700] <= 16'h0000;
      coeffs_in_data_log_force[ 701] <= 16'h0000;
      coeffs_in_data_log_force[ 702] <= 16'h0000;
      coeffs_in_data_log_force[ 703] <= 16'h0000;
      coeffs_in_data_log_force[ 704] <= 16'h0000;
      coeffs_in_data_log_force[ 705] <= 16'h0000;
      coeffs_in_data_log_force[ 706] <= 16'h0000;
      coeffs_in_data_log_force[ 707] <= 16'h0000;
      coeffs_in_data_log_force[ 708] <= 16'h0000;
      coeffs_in_data_log_force[ 709] <= 16'h0000;
      coeffs_in_data_log_force[ 710] <= 16'h0000;
      coeffs_in_data_log_force[ 711] <= 16'h0000;
      coeffs_in_data_log_force[ 712] <= 16'h0000;
      coeffs_in_data_log_force[ 713] <= 16'h0000;
      coeffs_in_data_log_force[ 714] <= 16'h0000;
      coeffs_in_data_log_force[ 715] <= 16'h0000;
      coeffs_in_data_log_force[ 716] <= 16'h0000;
      coeffs_in_data_log_force[ 717] <= 16'h0000;
      coeffs_in_data_log_force[ 718] <= 16'h0000;
      coeffs_in_data_log_force[ 719] <= 16'h0000;
      coeffs_in_data_log_force[ 720] <= 16'h0000;
      coeffs_in_data_log_force[ 721] <= 16'h0000;
      coeffs_in_data_log_force[ 722] <= 16'h0000;
      coeffs_in_data_log_force[ 723] <= 16'h0000;
      coeffs_in_data_log_force[ 724] <= 16'h0000;
      coeffs_in_data_log_force[ 725] <= 16'h0000;
      coeffs_in_data_log_force[ 726] <= 16'h0000;
      coeffs_in_data_log_force[ 727] <= 16'h0000;
      coeffs_in_data_log_force[ 728] <= 16'h0000;
      coeffs_in_data_log_force[ 729] <= 16'h0000;
      coeffs_in_data_log_force[ 730] <= 16'h0000;
      coeffs_in_data_log_force[ 731] <= 16'h0000;
      coeffs_in_data_log_force[ 732] <= 16'h0000;
      coeffs_in_data_log_force[ 733] <= 16'h0000;
      coeffs_in_data_log_force[ 734] <= 16'h0000;
      coeffs_in_data_log_force[ 735] <= 16'h0000;
      coeffs_in_data_log_force[ 736] <= 16'h0000;
      coeffs_in_data_log_force[ 737] <= 16'h0000;
      coeffs_in_data_log_force[ 738] <= 16'h0000;
      coeffs_in_data_log_force[ 739] <= 16'h0000;
      coeffs_in_data_log_force[ 740] <= 16'h0000;
      coeffs_in_data_log_force[ 741] <= 16'h0000;
      coeffs_in_data_log_force[ 742] <= 16'h0000;
      coeffs_in_data_log_force[ 743] <= 16'h0000;
      coeffs_in_data_log_force[ 744] <= 16'h0000;
      coeffs_in_data_log_force[ 745] <= 16'h0000;
      coeffs_in_data_log_force[ 746] <= 16'h0000;
      coeffs_in_data_log_force[ 747] <= 16'h0000;
      coeffs_in_data_log_force[ 748] <= 16'h0000;
      coeffs_in_data_log_force[ 749] <= 16'h0000;
      coeffs_in_data_log_force[ 750] <= 16'h0000;
      coeffs_in_data_log_force[ 751] <= 16'h0000;
      coeffs_in_data_log_force[ 752] <= 16'h0000;
      coeffs_in_data_log_force[ 753] <= 16'h0000;
      coeffs_in_data_log_force[ 754] <= 16'h0000;
      coeffs_in_data_log_force[ 755] <= 16'h0000;
      coeffs_in_data_log_force[ 756] <= 16'h0000;
      coeffs_in_data_log_force[ 757] <= 16'h0000;
      coeffs_in_data_log_force[ 758] <= 16'h0000;
      coeffs_in_data_log_force[ 759] <= 16'h0000;
      coeffs_in_data_log_force[ 760] <= 16'h0000;
      coeffs_in_data_log_force[ 761] <= 16'h0000;
      coeffs_in_data_log_force[ 762] <= 16'h0000;
      coeffs_in_data_log_force[ 763] <= 16'h0000;
      coeffs_in_data_log_force[ 764] <= 16'h0000;
      coeffs_in_data_log_force[ 765] <= 16'h0000;
      coeffs_in_data_log_force[ 766] <= 16'h0000;
      coeffs_in_data_log_force[ 767] <= 16'h0000;
      coeffs_in_data_log_force[ 768] <= 16'h0000;
      coeffs_in_data_log_force[ 769] <= 16'h0000;
      coeffs_in_data_log_force[ 770] <= 16'h0000;
      coeffs_in_data_log_force[ 771] <= 16'h0000;
      coeffs_in_data_log_force[ 772] <= 16'h0000;
      coeffs_in_data_log_force[ 773] <= 16'h0000;
      coeffs_in_data_log_force[ 774] <= 16'h0000;
      coeffs_in_data_log_force[ 775] <= 16'h0000;
      coeffs_in_data_log_force[ 776] <= 16'h0000;
      coeffs_in_data_log_force[ 777] <= 16'h0000;
      coeffs_in_data_log_force[ 778] <= 16'h0000;
      coeffs_in_data_log_force[ 779] <= 16'h0000;
      coeffs_in_data_log_force[ 780] <= 16'h0000;
      coeffs_in_data_log_force[ 781] <= 16'h0000;
      coeffs_in_data_log_force[ 782] <= 16'h0000;
      coeffs_in_data_log_force[ 783] <= 16'h0000;
      coeffs_in_data_log_force[ 784] <= 16'h0000;
      coeffs_in_data_log_force[ 785] <= 16'h0000;
      coeffs_in_data_log_force[ 786] <= 16'h0000;
      coeffs_in_data_log_force[ 787] <= 16'h0000;
      coeffs_in_data_log_force[ 788] <= 16'h0000;
      coeffs_in_data_log_force[ 789] <= 16'h0000;
      coeffs_in_data_log_force[ 790] <= 16'h0000;
      coeffs_in_data_log_force[ 791] <= 16'h0000;
      coeffs_in_data_log_force[ 792] <= 16'h0000;
      coeffs_in_data_log_force[ 793] <= 16'h0000;
      coeffs_in_data_log_force[ 794] <= 16'h0000;
      coeffs_in_data_log_force[ 795] <= 16'h0000;
      coeffs_in_data_log_force[ 796] <= 16'h0000;
      coeffs_in_data_log_force[ 797] <= 16'h0000;
      coeffs_in_data_log_force[ 798] <= 16'h0000;
      coeffs_in_data_log_force[ 799] <= 16'h0000;
      coeffs_in_data_log_force[ 800] <= 16'h0000;
      coeffs_in_data_log_force[ 801] <= 16'h0000;
      coeffs_in_data_log_force[ 802] <= 16'h0000;
      coeffs_in_data_log_force[ 803] <= 16'h0000;
      coeffs_in_data_log_force[ 804] <= 16'h0000;
      coeffs_in_data_log_force[ 805] <= 16'h0000;
      coeffs_in_data_log_force[ 806] <= 16'h0000;
      coeffs_in_data_log_force[ 807] <= 16'h0000;
      coeffs_in_data_log_force[ 808] <= 16'h0000;
      coeffs_in_data_log_force[ 809] <= 16'h0000;
      coeffs_in_data_log_force[ 810] <= 16'h0000;
      coeffs_in_data_log_force[ 811] <= 16'h0000;
      coeffs_in_data_log_force[ 812] <= 16'h0000;
      coeffs_in_data_log_force[ 813] <= 16'h0000;
      coeffs_in_data_log_force[ 814] <= 16'h0000;
      coeffs_in_data_log_force[ 815] <= 16'h0000;
      coeffs_in_data_log_force[ 816] <= 16'h0000;
      coeffs_in_data_log_force[ 817] <= 16'h0000;
      coeffs_in_data_log_force[ 818] <= 16'h0000;
      coeffs_in_data_log_force[ 819] <= 16'h0000;
      coeffs_in_data_log_force[ 820] <= 16'h0000;
      coeffs_in_data_log_force[ 821] <= 16'h0000;
      coeffs_in_data_log_force[ 822] <= 16'h0000;
      coeffs_in_data_log_force[ 823] <= 16'h0000;
      coeffs_in_data_log_force[ 824] <= 16'h0000;
      coeffs_in_data_log_force[ 825] <= 16'h0000;
      coeffs_in_data_log_force[ 826] <= 16'h0000;
      coeffs_in_data_log_force[ 827] <= 16'h0000;
      coeffs_in_data_log_force[ 828] <= 16'h0000;
      coeffs_in_data_log_force[ 829] <= 16'h0000;
      coeffs_in_data_log_force[ 830] <= 16'h0000;
      coeffs_in_data_log_force[ 831] <= 16'h0000;
      coeffs_in_data_log_force[ 832] <= 16'h0000;
      coeffs_in_data_log_force[ 833] <= 16'h0000;
      coeffs_in_data_log_force[ 834] <= 16'h0000;
      coeffs_in_data_log_force[ 835] <= 16'h0000;
      coeffs_in_data_log_force[ 836] <= 16'h0000;
      coeffs_in_data_log_force[ 837] <= 16'h0000;
      coeffs_in_data_log_force[ 838] <= 16'h0000;
      coeffs_in_data_log_force[ 839] <= 16'h0000;
      coeffs_in_data_log_force[ 840] <= 16'h0000;
      coeffs_in_data_log_force[ 841] <= 16'h0000;
      coeffs_in_data_log_force[ 842] <= 16'h0000;
      coeffs_in_data_log_force[ 843] <= 16'h0000;
      coeffs_in_data_log_force[ 844] <= 16'h0000;
      coeffs_in_data_log_force[ 845] <= 16'h0000;
      coeffs_in_data_log_force[ 846] <= 16'h0000;
      coeffs_in_data_log_force[ 847] <= 16'h0000;
      coeffs_in_data_log_force[ 848] <= 16'h0000;
      coeffs_in_data_log_force[ 849] <= 16'h0000;
      coeffs_in_data_log_force[ 850] <= 16'h0000;
      coeffs_in_data_log_force[ 851] <= 16'h0000;
      coeffs_in_data_log_force[ 852] <= 16'h0000;
      coeffs_in_data_log_force[ 853] <= 16'h0000;
      coeffs_in_data_log_force[ 854] <= 16'h0000;
      coeffs_in_data_log_force[ 855] <= 16'h0000;
      coeffs_in_data_log_force[ 856] <= 16'h0000;
      coeffs_in_data_log_force[ 857] <= 16'h0000;
      coeffs_in_data_log_force[ 858] <= 16'h0000;
      coeffs_in_data_log_force[ 859] <= 16'h0000;
      coeffs_in_data_log_force[ 860] <= 16'h0000;
      coeffs_in_data_log_force[ 861] <= 16'h0000;
      coeffs_in_data_log_force[ 862] <= 16'h0000;
      coeffs_in_data_log_force[ 863] <= 16'h0000;
      coeffs_in_data_log_force[ 864] <= 16'h0000;
      coeffs_in_data_log_force[ 865] <= 16'h0000;
      coeffs_in_data_log_force[ 866] <= 16'h0000;
      coeffs_in_data_log_force[ 867] <= 16'h0000;
      coeffs_in_data_log_force[ 868] <= 16'h0000;
      coeffs_in_data_log_force[ 869] <= 16'h0000;
      coeffs_in_data_log_force[ 870] <= 16'h0000;
      coeffs_in_data_log_force[ 871] <= 16'h0000;
      coeffs_in_data_log_force[ 872] <= 16'h0000;
      coeffs_in_data_log_force[ 873] <= 16'h0000;
      coeffs_in_data_log_force[ 874] <= 16'h0000;
      coeffs_in_data_log_force[ 875] <= 16'h0000;
      coeffs_in_data_log_force[ 876] <= 16'h0000;
      coeffs_in_data_log_force[ 877] <= 16'h0000;
      coeffs_in_data_log_force[ 878] <= 16'h0000;
      coeffs_in_data_log_force[ 879] <= 16'h0000;
      coeffs_in_data_log_force[ 880] <= 16'h0000;
      coeffs_in_data_log_force[ 881] <= 16'h0000;
      coeffs_in_data_log_force[ 882] <= 16'h0000;
      coeffs_in_data_log_force[ 883] <= 16'h0000;
      coeffs_in_data_log_force[ 884] <= 16'h0000;
      coeffs_in_data_log_force[ 885] <= 16'h0000;
      coeffs_in_data_log_force[ 886] <= 16'h0000;
      coeffs_in_data_log_force[ 887] <= 16'h0000;
      coeffs_in_data_log_force[ 888] <= 16'h0000;
      coeffs_in_data_log_force[ 889] <= 16'h0000;
      coeffs_in_data_log_force[ 890] <= 16'h0000;
      coeffs_in_data_log_force[ 891] <= 16'h0000;
      coeffs_in_data_log_force[ 892] <= 16'h0000;
      coeffs_in_data_log_force[ 893] <= 16'h0000;
      coeffs_in_data_log_force[ 894] <= 16'h0000;
      coeffs_in_data_log_force[ 895] <= 16'h0000;
      coeffs_in_data_log_force[ 896] <= 16'h0000;
      coeffs_in_data_log_force[ 897] <= 16'h0000;
      coeffs_in_data_log_force[ 898] <= 16'h0000;
      coeffs_in_data_log_force[ 899] <= 16'h0000;
      coeffs_in_data_log_force[ 900] <= 16'h0000;
      coeffs_in_data_log_force[ 901] <= 16'h0000;
      coeffs_in_data_log_force[ 902] <= 16'h0000;
      coeffs_in_data_log_force[ 903] <= 16'h0000;
      coeffs_in_data_log_force[ 904] <= 16'h0000;
      coeffs_in_data_log_force[ 905] <= 16'h0000;
      coeffs_in_data_log_force[ 906] <= 16'h0000;
      coeffs_in_data_log_force[ 907] <= 16'h0000;
      coeffs_in_data_log_force[ 908] <= 16'h0000;
      coeffs_in_data_log_force[ 909] <= 16'h0000;
      coeffs_in_data_log_force[ 910] <= 16'h0000;
      coeffs_in_data_log_force[ 911] <= 16'h0000;
      coeffs_in_data_log_force[ 912] <= 16'h0000;
      coeffs_in_data_log_force[ 913] <= 16'h0000;
      coeffs_in_data_log_force[ 914] <= 16'h0000;
      coeffs_in_data_log_force[ 915] <= 16'h0000;
      coeffs_in_data_log_force[ 916] <= 16'h0000;
      coeffs_in_data_log_force[ 917] <= 16'h0000;
      coeffs_in_data_log_force[ 918] <= 16'h0000;
      coeffs_in_data_log_force[ 919] <= 16'h0000;
      coeffs_in_data_log_force[ 920] <= 16'h0000;
      coeffs_in_data_log_force[ 921] <= 16'h0000;
      coeffs_in_data_log_force[ 922] <= 16'h0000;
      coeffs_in_data_log_force[ 923] <= 16'h0000;
      coeffs_in_data_log_force[ 924] <= 16'h0000;
      coeffs_in_data_log_force[ 925] <= 16'h0000;
      coeffs_in_data_log_force[ 926] <= 16'h0000;
      coeffs_in_data_log_force[ 927] <= 16'h0000;
      coeffs_in_data_log_force[ 928] <= 16'h0000;
      coeffs_in_data_log_force[ 929] <= 16'h0000;
      coeffs_in_data_log_force[ 930] <= 16'h0000;
      coeffs_in_data_log_force[ 931] <= 16'h0000;
      coeffs_in_data_log_force[ 932] <= 16'h0000;
      coeffs_in_data_log_force[ 933] <= 16'h0000;
      coeffs_in_data_log_force[ 934] <= 16'h0000;
      coeffs_in_data_log_force[ 935] <= 16'h0000;
      coeffs_in_data_log_force[ 936] <= 16'h0000;
      coeffs_in_data_log_force[ 937] <= 16'h0000;
      coeffs_in_data_log_force[ 938] <= 16'h0000;
      coeffs_in_data_log_force[ 939] <= 16'h0000;
      coeffs_in_data_log_force[ 940] <= 16'h0000;
      coeffs_in_data_log_force[ 941] <= 16'h0000;
      coeffs_in_data_log_force[ 942] <= 16'h0000;
      coeffs_in_data_log_force[ 943] <= 16'h0000;
      coeffs_in_data_log_force[ 944] <= 16'h0000;
      coeffs_in_data_log_force[ 945] <= 16'h0000;
      coeffs_in_data_log_force[ 946] <= 16'h0000;
      coeffs_in_data_log_force[ 947] <= 16'h0000;
      coeffs_in_data_log_force[ 948] <= 16'h0000;
      coeffs_in_data_log_force[ 949] <= 16'h0000;
      coeffs_in_data_log_force[ 950] <= 16'h0000;
      coeffs_in_data_log_force[ 951] <= 16'h0000;
      coeffs_in_data_log_force[ 952] <= 16'h0000;
      coeffs_in_data_log_force[ 953] <= 16'h0000;
      coeffs_in_data_log_force[ 954] <= 16'h0000;
      coeffs_in_data_log_force[ 955] <= 16'h0000;
      coeffs_in_data_log_force[ 956] <= 16'h0000;
      coeffs_in_data_log_force[ 957] <= 16'h0000;
      coeffs_in_data_log_force[ 958] <= 16'h0000;
      coeffs_in_data_log_force[ 959] <= 16'h0000;
      coeffs_in_data_log_force[ 960] <= 16'h0000;
      coeffs_in_data_log_force[ 961] <= 16'h0000;
      coeffs_in_data_log_force[ 962] <= 16'h0000;
      coeffs_in_data_log_force[ 963] <= 16'h0000;
      coeffs_in_data_log_force[ 964] <= 16'h0000;
      coeffs_in_data_log_force[ 965] <= 16'h0000;
      coeffs_in_data_log_force[ 966] <= 16'h0000;
      coeffs_in_data_log_force[ 967] <= 16'h0000;
      coeffs_in_data_log_force[ 968] <= 16'h0000;
      coeffs_in_data_log_force[ 969] <= 16'h0000;
      coeffs_in_data_log_force[ 970] <= 16'h0000;
      coeffs_in_data_log_force[ 971] <= 16'h0000;
      coeffs_in_data_log_force[ 972] <= 16'h0000;
      coeffs_in_data_log_force[ 973] <= 16'h0000;
      coeffs_in_data_log_force[ 974] <= 16'h0000;
      coeffs_in_data_log_force[ 975] <= 16'h0000;
      coeffs_in_data_log_force[ 976] <= 16'h0000;
      coeffs_in_data_log_force[ 977] <= 16'h0000;
      coeffs_in_data_log_force[ 978] <= 16'h0000;
      coeffs_in_data_log_force[ 979] <= 16'h0000;
      coeffs_in_data_log_force[ 980] <= 16'h0000;
      coeffs_in_data_log_force[ 981] <= 16'h0000;
      coeffs_in_data_log_force[ 982] <= 16'h0000;
      coeffs_in_data_log_force[ 983] <= 16'h0000;
      coeffs_in_data_log_force[ 984] <= 16'h0000;
      coeffs_in_data_log_force[ 985] <= 16'h0000;
      coeffs_in_data_log_force[ 986] <= 16'h0000;
      coeffs_in_data_log_force[ 987] <= 16'h0000;
      coeffs_in_data_log_force[ 988] <= 16'h0000;
      coeffs_in_data_log_force[ 989] <= 16'h0000;
      coeffs_in_data_log_force[ 990] <= 16'h0000;
      coeffs_in_data_log_force[ 991] <= 16'h0000;
      coeffs_in_data_log_force[ 992] <= 16'h0000;
      coeffs_in_data_log_force[ 993] <= 16'h0000;
      coeffs_in_data_log_force[ 994] <= 16'h0000;
      coeffs_in_data_log_force[ 995] <= 16'h0000;
      coeffs_in_data_log_force[ 996] <= 16'h0000;
      coeffs_in_data_log_force[ 997] <= 16'h0000;
      coeffs_in_data_log_force[ 998] <= 16'h0000;
      coeffs_in_data_log_force[ 999] <= 16'h0000;
      coeffs_in_data_log_force[1000] <= 16'h0000;
      coeffs_in_data_log_force[1001] <= 16'h0000;
      coeffs_in_data_log_force[1002] <= 16'h0000;
      coeffs_in_data_log_force[1003] <= 16'h0000;
      coeffs_in_data_log_force[1004] <= 16'h0000;
      coeffs_in_data_log_force[1005] <= 16'h0000;
      coeffs_in_data_log_force[1006] <= 16'h0000;
      coeffs_in_data_log_force[1007] <= 16'h0000;
      coeffs_in_data_log_force[1008] <= 16'h0000;
      coeffs_in_data_log_force[1009] <= 16'h0000;
      coeffs_in_data_log_force[1010] <= 16'h0000;
      coeffs_in_data_log_force[1011] <= 16'h0000;
      coeffs_in_data_log_force[1012] <= 16'h0000;
      coeffs_in_data_log_force[1013] <= 16'h0000;
      coeffs_in_data_log_force[1014] <= 16'h0000;
      coeffs_in_data_log_force[1015] <= 16'h0000;
      coeffs_in_data_log_force[1016] <= 16'h0000;
      coeffs_in_data_log_force[1017] <= 16'h0000;
      coeffs_in_data_log_force[1018] <= 16'h0000;
      coeffs_in_data_log_force[1019] <= 16'h0000;
      coeffs_in_data_log_force[1020] <= 16'h0000;
      coeffs_in_data_log_force[1021] <= 16'h0000;
      coeffs_in_data_log_force[1022] <= 16'h0000;
      coeffs_in_data_log_force[1023] <= 16'h0000;
      coeffs_in_data_log_force[1024] <= 16'h0000;
      coeffs_in_data_log_force[1025] <= 16'h0000;
      coeffs_in_data_log_force[1026] <= 16'h0000;
      coeffs_in_data_log_force[1027] <= 16'h0000;
      coeffs_in_data_log_force[1028] <= 16'h0000;
      coeffs_in_data_log_force[1029] <= 16'h0000;
      coeffs_in_data_log_force[1030] <= 16'h0000;
      coeffs_in_data_log_force[1031] <= 16'h0000;
      coeffs_in_data_log_force[1032] <= 16'h0000;
      coeffs_in_data_log_force[1033] <= 16'h0000;
      coeffs_in_data_log_force[1034] <= 16'h0000;
      coeffs_in_data_log_force[1035] <= 16'h0000;
      coeffs_in_data_log_force[1036] <= 16'h0000;
      coeffs_in_data_log_force[1037] <= 16'h0000;
      coeffs_in_data_log_force[1038] <= 16'h0000;
      coeffs_in_data_log_force[1039] <= 16'h0000;
      coeffs_in_data_log_force[1040] <= 16'h0000;
      coeffs_in_data_log_force[1041] <= 16'h0000;
      coeffs_in_data_log_force[1042] <= 16'h0000;
      coeffs_in_data_log_force[1043] <= 16'h0000;
      coeffs_in_data_log_force[1044] <= 16'h0000;
      coeffs_in_data_log_force[1045] <= 16'h0000;
      coeffs_in_data_log_force[1046] <= 16'h0000;
      coeffs_in_data_log_force[1047] <= 16'h0000;
      coeffs_in_data_log_force[1048] <= 16'h0000;
      coeffs_in_data_log_force[1049] <= 16'h0000;
      coeffs_in_data_log_force[1050] <= 16'h0000;
      coeffs_in_data_log_force[1051] <= 16'h0000;
      coeffs_in_data_log_force[1052] <= 16'h0000;
      coeffs_in_data_log_force[1053] <= 16'h0000;
      coeffs_in_data_log_force[1054] <= 16'h0000;
      coeffs_in_data_log_force[1055] <= 16'h0000;
      coeffs_in_data_log_force[1056] <= 16'h0000;
      coeffs_in_data_log_force[1057] <= 16'h0000;
      coeffs_in_data_log_force[1058] <= 16'h0000;
      coeffs_in_data_log_force[1059] <= 16'h0000;
      coeffs_in_data_log_force[1060] <= 16'h0000;
      coeffs_in_data_log_force[1061] <= 16'h0000;
      coeffs_in_data_log_force[1062] <= 16'h0000;
      coeffs_in_data_log_force[1063] <= 16'h0000;
      coeffs_in_data_log_force[1064] <= 16'h0000;
      coeffs_in_data_log_force[1065] <= 16'h0000;
      coeffs_in_data_log_force[1066] <= 16'h0000;
      coeffs_in_data_log_force[1067] <= 16'h0000;
      coeffs_in_data_log_force[1068] <= 16'h0000;
      coeffs_in_data_log_force[1069] <= 16'h0000;
      coeffs_in_data_log_force[1070] <= 16'h0000;
      coeffs_in_data_log_force[1071] <= 16'h0000;
      coeffs_in_data_log_force[1072] <= 16'h0000;
      coeffs_in_data_log_force[1073] <= 16'h0000;
      coeffs_in_data_log_force[1074] <= 16'h0000;
      coeffs_in_data_log_force[1075] <= 16'h0000;
      coeffs_in_data_log_force[1076] <= 16'h0000;
      coeffs_in_data_log_force[1077] <= 16'h0000;
      coeffs_in_data_log_force[1078] <= 16'h0000;
      coeffs_in_data_log_force[1079] <= 16'h0000;
      coeffs_in_data_log_force[1080] <= 16'h0000;
      coeffs_in_data_log_force[1081] <= 16'h0000;
      coeffs_in_data_log_force[1082] <= 16'h0000;
      coeffs_in_data_log_force[1083] <= 16'h0000;
      coeffs_in_data_log_force[1084] <= 16'h0000;
      coeffs_in_data_log_force[1085] <= 16'h0000;
      coeffs_in_data_log_force[1086] <= 16'h0000;
      coeffs_in_data_log_force[1087] <= 16'h0000;
      coeffs_in_data_log_force[1088] <= 16'h0000;
      coeffs_in_data_log_force[1089] <= 16'h0000;
      coeffs_in_data_log_force[1090] <= 16'h0000;
      coeffs_in_data_log_force[1091] <= 16'h0000;
      coeffs_in_data_log_force[1092] <= 16'h0000;
      coeffs_in_data_log_force[1093] <= 16'h0000;
      coeffs_in_data_log_force[1094] <= 16'h0000;
      coeffs_in_data_log_force[1095] <= 16'h0000;
      coeffs_in_data_log_force[1096] <= 16'h0000;
      coeffs_in_data_log_force[1097] <= 16'h0000;
      coeffs_in_data_log_force[1098] <= 16'h0000;
      coeffs_in_data_log_force[1099] <= 16'h0000;
      coeffs_in_data_log_force[1100] <= 16'h0000;
      coeffs_in_data_log_force[1101] <= 16'h0000;
      coeffs_in_data_log_force[1102] <= 16'h0000;
      coeffs_in_data_log_force[1103] <= 16'h0000;
      coeffs_in_data_log_force[1104] <= 16'h0000;
      coeffs_in_data_log_force[1105] <= 16'h0000;
      coeffs_in_data_log_force[1106] <= 16'h0000;
      coeffs_in_data_log_force[1107] <= 16'h0000;
      coeffs_in_data_log_force[1108] <= 16'h0000;
      coeffs_in_data_log_force[1109] <= 16'h0000;
      coeffs_in_data_log_force[1110] <= 16'h0000;
      coeffs_in_data_log_force[1111] <= 16'h0000;
      coeffs_in_data_log_force[1112] <= 16'h0000;
      coeffs_in_data_log_force[1113] <= 16'h0000;
      coeffs_in_data_log_force[1114] <= 16'h0000;
      coeffs_in_data_log_force[1115] <= 16'h0000;
      coeffs_in_data_log_force[1116] <= 16'h0000;
      coeffs_in_data_log_force[1117] <= 16'h0000;
      coeffs_in_data_log_force[1118] <= 16'h0000;
      coeffs_in_data_log_force[1119] <= 16'h0000;
      coeffs_in_data_log_force[1120] <= 16'h0000;
      coeffs_in_data_log_force[1121] <= 16'h0000;
      coeffs_in_data_log_force[1122] <= 16'h0000;
      coeffs_in_data_log_force[1123] <= 16'h0000;
      coeffs_in_data_log_force[1124] <= 16'h0000;
      coeffs_in_data_log_force[1125] <= 16'h0000;
      coeffs_in_data_log_force[1126] <= 16'h0000;
      coeffs_in_data_log_force[1127] <= 16'h0000;
      coeffs_in_data_log_force[1128] <= 16'h0000;
      coeffs_in_data_log_force[1129] <= 16'h0000;
      coeffs_in_data_log_force[1130] <= 16'h0000;
      coeffs_in_data_log_force[1131] <= 16'h0000;
      coeffs_in_data_log_force[1132] <= 16'h0000;
      coeffs_in_data_log_force[1133] <= 16'h0000;
      coeffs_in_data_log_force[1134] <= 16'h0000;
      coeffs_in_data_log_force[1135] <= 16'h0000;
      coeffs_in_data_log_force[1136] <= 16'h0000;
      coeffs_in_data_log_force[1137] <= 16'h0000;
      coeffs_in_data_log_force[1138] <= 16'h0000;
      coeffs_in_data_log_force[1139] <= 16'h0000;
      coeffs_in_data_log_force[1140] <= 16'h0000;
      coeffs_in_data_log_force[1141] <= 16'h0000;
      coeffs_in_data_log_force[1142] <= 16'h0000;
      coeffs_in_data_log_force[1143] <= 16'h0000;
      coeffs_in_data_log_force[1144] <= 16'h0000;
      coeffs_in_data_log_force[1145] <= 16'h0000;
      coeffs_in_data_log_force[1146] <= 16'h0000;
      coeffs_in_data_log_force[1147] <= 16'h0000;
      coeffs_in_data_log_force[1148] <= 16'h0000;
      coeffs_in_data_log_force[1149] <= 16'h0000;
      coeffs_in_data_log_force[1150] <= 16'h0000;
      coeffs_in_data_log_force[1151] <= 16'h0000;
      coeffs_in_data_log_force[1152] <= 16'h0000;
      coeffs_in_data_log_force[1153] <= 16'h0000;
      coeffs_in_data_log_force[1154] <= 16'h0000;
      coeffs_in_data_log_force[1155] <= 16'h0000;
      coeffs_in_data_log_force[1156] <= 16'h0000;
      coeffs_in_data_log_force[1157] <= 16'h0000;
      coeffs_in_data_log_force[1158] <= 16'h0000;
      coeffs_in_data_log_force[1159] <= 16'h0000;
      coeffs_in_data_log_force[1160] <= 16'h0000;
      coeffs_in_data_log_force[1161] <= 16'h0000;
      coeffs_in_data_log_force[1162] <= 16'h0000;
      coeffs_in_data_log_force[1163] <= 16'h0000;
      coeffs_in_data_log_force[1164] <= 16'h0000;
      coeffs_in_data_log_force[1165] <= 16'h0000;
      coeffs_in_data_log_force[1166] <= 16'h0000;
      coeffs_in_data_log_force[1167] <= 16'h0000;
      coeffs_in_data_log_force[1168] <= 16'h0000;
      coeffs_in_data_log_force[1169] <= 16'h0000;
      coeffs_in_data_log_force[1170] <= 16'h0000;
      coeffs_in_data_log_force[1171] <= 16'h0000;
      coeffs_in_data_log_force[1172] <= 16'h0000;
      coeffs_in_data_log_force[1173] <= 16'h0000;
      coeffs_in_data_log_force[1174] <= 16'h0000;
      coeffs_in_data_log_force[1175] <= 16'h0000;
      coeffs_in_data_log_force[1176] <= 16'h0000;
      coeffs_in_data_log_force[1177] <= 16'h0000;
      coeffs_in_data_log_force[1178] <= 16'h0000;
      coeffs_in_data_log_force[1179] <= 16'h0000;
      coeffs_in_data_log_force[1180] <= 16'h0000;
      coeffs_in_data_log_force[1181] <= 16'h0000;
      coeffs_in_data_log_force[1182] <= 16'h0000;
      coeffs_in_data_log_force[1183] <= 16'h0000;
      coeffs_in_data_log_force[1184] <= 16'h0000;
      coeffs_in_data_log_force[1185] <= 16'h0000;
      coeffs_in_data_log_force[1186] <= 16'h0000;
      coeffs_in_data_log_force[1187] <= 16'h0000;
      coeffs_in_data_log_force[1188] <= 16'h0000;
      coeffs_in_data_log_force[1189] <= 16'h0000;
      coeffs_in_data_log_force[1190] <= 16'h0000;
      coeffs_in_data_log_force[1191] <= 16'h0000;
      coeffs_in_data_log_force[1192] <= 16'h0000;
      coeffs_in_data_log_force[1193] <= 16'h0000;
      coeffs_in_data_log_force[1194] <= 16'h0000;
      coeffs_in_data_log_force[1195] <= 16'h0000;
      coeffs_in_data_log_force[1196] <= 16'h0000;
      coeffs_in_data_log_force[1197] <= 16'h0000;
      coeffs_in_data_log_force[1198] <= 16'h0000;
      coeffs_in_data_log_force[1199] <= 16'h0000;
      coeffs_in_data_log_force[1200] <= 16'h0000;
      coeffs_in_data_log_force[1201] <= 16'h0000;
      coeffs_in_data_log_force[1202] <= 16'h0000;
      coeffs_in_data_log_force[1203] <= 16'h0000;
      coeffs_in_data_log_force[1204] <= 16'h0000;
      coeffs_in_data_log_force[1205] <= 16'h0000;
      coeffs_in_data_log_force[1206] <= 16'h0000;
      coeffs_in_data_log_force[1207] <= 16'h0000;
      coeffs_in_data_log_force[1208] <= 16'h0000;
      coeffs_in_data_log_force[1209] <= 16'h0000;
      coeffs_in_data_log_force[1210] <= 16'h0000;
      coeffs_in_data_log_force[1211] <= 16'h0000;
      coeffs_in_data_log_force[1212] <= 16'h0000;
      coeffs_in_data_log_force[1213] <= 16'h0000;
      coeffs_in_data_log_force[1214] <= 16'h0000;
      coeffs_in_data_log_force[1215] <= 16'h0000;
      coeffs_in_data_log_force[1216] <= 16'h0000;
      coeffs_in_data_log_force[1217] <= 16'h0000;
      coeffs_in_data_log_force[1218] <= 16'h0000;
      coeffs_in_data_log_force[1219] <= 16'h0000;
      coeffs_in_data_log_force[1220] <= 16'h0000;
      coeffs_in_data_log_force[1221] <= 16'h0000;
      coeffs_in_data_log_force[1222] <= 16'h0000;
      coeffs_in_data_log_force[1223] <= 16'h0000;
      coeffs_in_data_log_force[1224] <= 16'h0000;
      coeffs_in_data_log_force[1225] <= 16'h0000;
      coeffs_in_data_log_force[1226] <= 16'h0000;
      coeffs_in_data_log_force[1227] <= 16'h0000;
      coeffs_in_data_log_force[1228] <= 16'h0000;
      coeffs_in_data_log_force[1229] <= 16'h0000;
      coeffs_in_data_log_force[1230] <= 16'h0000;
      coeffs_in_data_log_force[1231] <= 16'h0000;
      coeffs_in_data_log_force[1232] <= 16'h0000;
      coeffs_in_data_log_force[1233] <= 16'h0000;
      coeffs_in_data_log_force[1234] <= 16'h0000;
      coeffs_in_data_log_force[1235] <= 16'h0000;
      coeffs_in_data_log_force[1236] <= 16'h0000;
      coeffs_in_data_log_force[1237] <= 16'h0000;
      coeffs_in_data_log_force[1238] <= 16'h0000;
      coeffs_in_data_log_force[1239] <= 16'h0000;
      coeffs_in_data_log_force[1240] <= 16'h0000;
      coeffs_in_data_log_force[1241] <= 16'h0000;
      coeffs_in_data_log_force[1242] <= 16'h0000;
      coeffs_in_data_log_force[1243] <= 16'h0000;
      coeffs_in_data_log_force[1244] <= 16'h0000;
      coeffs_in_data_log_force[1245] <= 16'h0000;
      coeffs_in_data_log_force[1246] <= 16'h0000;
      coeffs_in_data_log_force[1247] <= 16'h0000;
      coeffs_in_data_log_force[1248] <= 16'h0000;
      coeffs_in_data_log_force[1249] <= 16'h0000;
      coeffs_in_data_log_force[1250] <= 16'h0000;
      coeffs_in_data_log_force[1251] <= 16'h0000;
      coeffs_in_data_log_force[1252] <= 16'h0000;
      coeffs_in_data_log_force[1253] <= 16'h0000;
      coeffs_in_data_log_force[1254] <= 16'h0000;
      coeffs_in_data_log_force[1255] <= 16'h0000;
      coeffs_in_data_log_force[1256] <= 16'h0000;
      coeffs_in_data_log_force[1257] <= 16'h0000;
      coeffs_in_data_log_force[1258] <= 16'h0000;
      coeffs_in_data_log_force[1259] <= 16'h0000;
      coeffs_in_data_log_force[1260] <= 16'h0000;
      coeffs_in_data_log_force[1261] <= 16'h0000;
      coeffs_in_data_log_force[1262] <= 16'h0000;
      coeffs_in_data_log_force[1263] <= 16'h0000;
      coeffs_in_data_log_force[1264] <= 16'h0000;
      coeffs_in_data_log_force[1265] <= 16'h0000;
      coeffs_in_data_log_force[1266] <= 16'h0000;
      coeffs_in_data_log_force[1267] <= 16'h0000;
      coeffs_in_data_log_force[1268] <= 16'h0000;
      coeffs_in_data_log_force[1269] <= 16'h0000;
      coeffs_in_data_log_force[1270] <= 16'h0000;
      coeffs_in_data_log_force[1271] <= 16'h0000;
      coeffs_in_data_log_force[1272] <= 16'h0000;
      coeffs_in_data_log_force[1273] <= 16'h0000;
      coeffs_in_data_log_force[1274] <= 16'h0000;
      coeffs_in_data_log_force[1275] <= 16'h0000;
      coeffs_in_data_log_force[1276] <= 16'h0000;
      coeffs_in_data_log_force[1277] <= 16'h0000;
      coeffs_in_data_log_force[1278] <= 16'h0000;
      coeffs_in_data_log_force[1279] <= 16'h0000;
      coeffs_in_data_log_force[1280] <= 16'h0000;
      coeffs_in_data_log_force[1281] <= 16'h0000;
      coeffs_in_data_log_force[1282] <= 16'h0000;
      coeffs_in_data_log_force[1283] <= 16'h0000;
      coeffs_in_data_log_force[1284] <= 16'h0000;
      coeffs_in_data_log_force[1285] <= 16'h0000;
      coeffs_in_data_log_force[1286] <= 16'h0000;
      coeffs_in_data_log_force[1287] <= 16'h0000;
      coeffs_in_data_log_force[1288] <= 16'h0000;
      coeffs_in_data_log_force[1289] <= 16'h0000;
      coeffs_in_data_log_force[1290] <= 16'h0000;
      coeffs_in_data_log_force[1291] <= 16'h0000;
      coeffs_in_data_log_force[1292] <= 16'h0000;
      coeffs_in_data_log_force[1293] <= 16'h0000;
      coeffs_in_data_log_force[1294] <= 16'h0000;
      coeffs_in_data_log_force[1295] <= 16'h0000;
      coeffs_in_data_log_force[1296] <= 16'h0000;
      coeffs_in_data_log_force[1297] <= 16'h0000;
      coeffs_in_data_log_force[1298] <= 16'h0000;
      coeffs_in_data_log_force[1299] <= 16'h0000;
      coeffs_in_data_log_force[1300] <= 16'h0000;
      coeffs_in_data_log_force[1301] <= 16'h0000;
      coeffs_in_data_log_force[1302] <= 16'h0000;
      coeffs_in_data_log_force[1303] <= 16'h0000;
      coeffs_in_data_log_force[1304] <= 16'h0000;
      coeffs_in_data_log_force[1305] <= 16'h0000;
      coeffs_in_data_log_force[1306] <= 16'h0000;
      coeffs_in_data_log_force[1307] <= 16'h0000;
      coeffs_in_data_log_force[1308] <= 16'h0000;
      coeffs_in_data_log_force[1309] <= 16'h0000;
      coeffs_in_data_log_force[1310] <= 16'h0000;
      coeffs_in_data_log_force[1311] <= 16'h0000;
      coeffs_in_data_log_force[1312] <= 16'h0000;
      coeffs_in_data_log_force[1313] <= 16'h0000;
      coeffs_in_data_log_force[1314] <= 16'h0000;
      coeffs_in_data_log_force[1315] <= 16'h0000;
      coeffs_in_data_log_force[1316] <= 16'h0000;
      coeffs_in_data_log_force[1317] <= 16'h0000;
      coeffs_in_data_log_force[1318] <= 16'h0000;
      coeffs_in_data_log_force[1319] <= 16'h0000;
      coeffs_in_data_log_force[1320] <= 16'h0000;
      coeffs_in_data_log_force[1321] <= 16'h0000;
      coeffs_in_data_log_force[1322] <= 16'h0000;
      coeffs_in_data_log_force[1323] <= 16'h0000;
      coeffs_in_data_log_force[1324] <= 16'h0000;
      coeffs_in_data_log_force[1325] <= 16'h0000;
      coeffs_in_data_log_force[1326] <= 16'h0000;
      coeffs_in_data_log_force[1327] <= 16'h0000;
      coeffs_in_data_log_force[1328] <= 16'h0000;
      coeffs_in_data_log_force[1329] <= 16'h0000;
      coeffs_in_data_log_force[1330] <= 16'h0000;
      coeffs_in_data_log_force[1331] <= 16'h0000;
      coeffs_in_data_log_force[1332] <= 16'h0000;
      coeffs_in_data_log_force[1333] <= 16'h0000;
      coeffs_in_data_log_force[1334] <= 16'h0000;
      coeffs_in_data_log_force[1335] <= 16'h0000;
      coeffs_in_data_log_force[1336] <= 16'h0000;
      coeffs_in_data_log_force[1337] <= 16'h0000;
      coeffs_in_data_log_force[1338] <= 16'h0000;
      coeffs_in_data_log_force[1339] <= 16'h0000;
      coeffs_in_data_log_force[1340] <= 16'h0000;
      coeffs_in_data_log_force[1341] <= 16'h0000;
      coeffs_in_data_log_force[1342] <= 16'h0000;
      coeffs_in_data_log_force[1343] <= 16'h0000;
      coeffs_in_data_log_force[1344] <= 16'h0000;
      coeffs_in_data_log_force[1345] <= 16'h0000;
      coeffs_in_data_log_force[1346] <= 16'h0000;
      coeffs_in_data_log_force[1347] <= 16'h0000;
      coeffs_in_data_log_force[1348] <= 16'h0000;
      coeffs_in_data_log_force[1349] <= 16'h0000;
      coeffs_in_data_log_force[1350] <= 16'h0000;
      coeffs_in_data_log_force[1351] <= 16'h0000;
      coeffs_in_data_log_force[1352] <= 16'h0000;
      coeffs_in_data_log_force[1353] <= 16'h0000;
      coeffs_in_data_log_force[1354] <= 16'h0000;
      coeffs_in_data_log_force[1355] <= 16'h0000;
      coeffs_in_data_log_force[1356] <= 16'h0000;
      coeffs_in_data_log_force[1357] <= 16'h0000;
      coeffs_in_data_log_force[1358] <= 16'h0000;
      coeffs_in_data_log_force[1359] <= 16'h0000;
      coeffs_in_data_log_force[1360] <= 16'h0000;
      coeffs_in_data_log_force[1361] <= 16'h0000;
      coeffs_in_data_log_force[1362] <= 16'h0000;
      coeffs_in_data_log_force[1363] <= 16'h0000;
      coeffs_in_data_log_force[1364] <= 16'h0000;
      coeffs_in_data_log_force[1365] <= 16'h0000;
      coeffs_in_data_log_force[1366] <= 16'h0000;
      coeffs_in_data_log_force[1367] <= 16'h0000;
      coeffs_in_data_log_force[1368] <= 16'h0000;
      coeffs_in_data_log_force[1369] <= 16'h0000;
      coeffs_in_data_log_force[1370] <= 16'h0000;
      coeffs_in_data_log_force[1371] <= 16'h0000;
      coeffs_in_data_log_force[1372] <= 16'h0000;
      coeffs_in_data_log_force[1373] <= 16'h0000;
      coeffs_in_data_log_force[1374] <= 16'h0000;
      coeffs_in_data_log_force[1375] <= 16'h0000;
      coeffs_in_data_log_force[1376] <= 16'h0000;
      coeffs_in_data_log_force[1377] <= 16'h0000;
      coeffs_in_data_log_force[1378] <= 16'h0000;
      coeffs_in_data_log_force[1379] <= 16'h0000;
      coeffs_in_data_log_force[1380] <= 16'h0000;
      coeffs_in_data_log_force[1381] <= 16'h0000;
      coeffs_in_data_log_force[1382] <= 16'h0000;
      coeffs_in_data_log_force[1383] <= 16'h0000;
      coeffs_in_data_log_force[1384] <= 16'h0000;
      coeffs_in_data_log_force[1385] <= 16'h0000;
      coeffs_in_data_log_force[1386] <= 16'h0000;
      coeffs_in_data_log_force[1387] <= 16'h0000;
      coeffs_in_data_log_force[1388] <= 16'h0000;
      coeffs_in_data_log_force[1389] <= 16'h0000;
      coeffs_in_data_log_force[1390] <= 16'h0000;
      coeffs_in_data_log_force[1391] <= 16'h0000;
      coeffs_in_data_log_force[1392] <= 16'h0000;
      coeffs_in_data_log_force[1393] <= 16'h0000;
      coeffs_in_data_log_force[1394] <= 16'h0000;
      coeffs_in_data_log_force[1395] <= 16'h0000;
      coeffs_in_data_log_force[1396] <= 16'h0000;
      coeffs_in_data_log_force[1397] <= 16'h0000;
      coeffs_in_data_log_force[1398] <= 16'h0000;
      coeffs_in_data_log_force[1399] <= 16'h0000;
      coeffs_in_data_log_force[1400] <= 16'h0000;
      coeffs_in_data_log_force[1401] <= 16'h0000;
      coeffs_in_data_log_force[1402] <= 16'h0000;
      coeffs_in_data_log_force[1403] <= 16'h0000;
      coeffs_in_data_log_force[1404] <= 16'h0000;
      coeffs_in_data_log_force[1405] <= 16'h0000;
      coeffs_in_data_log_force[1406] <= 16'h0000;
      coeffs_in_data_log_force[1407] <= 16'h0000;
      coeffs_in_data_log_force[1408] <= 16'h0000;
      coeffs_in_data_log_force[1409] <= 16'h0000;
      coeffs_in_data_log_force[1410] <= 16'h0000;
      coeffs_in_data_log_force[1411] <= 16'h0000;
      coeffs_in_data_log_force[1412] <= 16'h0000;
      coeffs_in_data_log_force[1413] <= 16'h0000;
      coeffs_in_data_log_force[1414] <= 16'h0000;
      coeffs_in_data_log_force[1415] <= 16'h0000;
      coeffs_in_data_log_force[1416] <= 16'h0000;
      coeffs_in_data_log_force[1417] <= 16'h0000;
      coeffs_in_data_log_force[1418] <= 16'h0000;
      coeffs_in_data_log_force[1419] <= 16'h0000;
      coeffs_in_data_log_force[1420] <= 16'h0000;
      coeffs_in_data_log_force[1421] <= 16'h0000;
      coeffs_in_data_log_force[1422] <= 16'h0000;
      coeffs_in_data_log_force[1423] <= 16'h0000;
      coeffs_in_data_log_force[1424] <= 16'h0000;
      coeffs_in_data_log_force[1425] <= 16'h0000;
      coeffs_in_data_log_force[1426] <= 16'h0000;
      coeffs_in_data_log_force[1427] <= 16'h0000;
      coeffs_in_data_log_force[1428] <= 16'h0000;
      coeffs_in_data_log_force[1429] <= 16'h0000;
      coeffs_in_data_log_force[1430] <= 16'h0000;
      coeffs_in_data_log_force[1431] <= 16'h0000;
      coeffs_in_data_log_force[1432] <= 16'h0000;
      coeffs_in_data_log_force[1433] <= 16'h0000;
      coeffs_in_data_log_force[1434] <= 16'h0000;
      coeffs_in_data_log_force[1435] <= 16'h0000;
      coeffs_in_data_log_force[1436] <= 16'h0000;
      coeffs_in_data_log_force[1437] <= 16'h0000;
      coeffs_in_data_log_force[1438] <= 16'h0000;
      coeffs_in_data_log_force[1439] <= 16'h0000;
      coeffs_in_data_log_force[1440] <= 16'h0000;
      coeffs_in_data_log_force[1441] <= 16'h0000;
      coeffs_in_data_log_force[1442] <= 16'h0000;
      coeffs_in_data_log_force[1443] <= 16'h0000;
      coeffs_in_data_log_force[1444] <= 16'h0000;
      coeffs_in_data_log_force[1445] <= 16'h0000;
      coeffs_in_data_log_force[1446] <= 16'h0000;
      coeffs_in_data_log_force[1447] <= 16'h0000;
      coeffs_in_data_log_force[1448] <= 16'h0000;
      coeffs_in_data_log_force[1449] <= 16'h0000;
      coeffs_in_data_log_force[1450] <= 16'h0000;
      coeffs_in_data_log_force[1451] <= 16'h0000;
      coeffs_in_data_log_force[1452] <= 16'h0000;
      coeffs_in_data_log_force[1453] <= 16'h0000;
      coeffs_in_data_log_force[1454] <= 16'h0000;
      coeffs_in_data_log_force[1455] <= 16'h0000;
      coeffs_in_data_log_force[1456] <= 16'h0000;
      coeffs_in_data_log_force[1457] <= 16'h0000;
      coeffs_in_data_log_force[1458] <= 16'h0000;
      coeffs_in_data_log_force[1459] <= 16'h0000;
      coeffs_in_data_log_force[1460] <= 16'h0000;
      coeffs_in_data_log_force[1461] <= 16'h0000;
      coeffs_in_data_log_force[1462] <= 16'h0000;
      coeffs_in_data_log_force[1463] <= 16'h0000;
      coeffs_in_data_log_force[1464] <= 16'h0000;
      coeffs_in_data_log_force[1465] <= 16'h0000;
      coeffs_in_data_log_force[1466] <= 16'h0000;
      coeffs_in_data_log_force[1467] <= 16'h0000;
      coeffs_in_data_log_force[1468] <= 16'h0000;
      coeffs_in_data_log_force[1469] <= 16'h0000;
      coeffs_in_data_log_force[1470] <= 16'h0000;
      coeffs_in_data_log_force[1471] <= 16'h0000;
      coeffs_in_data_log_force[1472] <= 16'h0000;
      coeffs_in_data_log_force[1473] <= 16'h0000;
      coeffs_in_data_log_force[1474] <= 16'h0000;
      coeffs_in_data_log_force[1475] <= 16'h0000;
      coeffs_in_data_log_force[1476] <= 16'h0000;
      coeffs_in_data_log_force[1477] <= 16'h0000;
      coeffs_in_data_log_force[1478] <= 16'h0000;
      coeffs_in_data_log_force[1479] <= 16'h0000;
      coeffs_in_data_log_force[1480] <= 16'h0000;
      coeffs_in_data_log_force[1481] <= 16'h0000;
      coeffs_in_data_log_force[1482] <= 16'h0000;
      coeffs_in_data_log_force[1483] <= 16'h0000;
      coeffs_in_data_log_force[1484] <= 16'h0000;
      coeffs_in_data_log_force[1485] <= 16'h0000;
      coeffs_in_data_log_force[1486] <= 16'h0000;
      coeffs_in_data_log_force[1487] <= 16'h0000;
      coeffs_in_data_log_force[1488] <= 16'h0000;
      coeffs_in_data_log_force[1489] <= 16'h0000;
      coeffs_in_data_log_force[1490] <= 16'h0000;
      coeffs_in_data_log_force[1491] <= 16'h0000;
      coeffs_in_data_log_force[1492] <= 16'h0000;
      coeffs_in_data_log_force[1493] <= 16'h0000;
      coeffs_in_data_log_force[1494] <= 16'h0000;
      coeffs_in_data_log_force[1495] <= 16'h0000;
      coeffs_in_data_log_force[1496] <= 16'h0000;
      coeffs_in_data_log_force[1497] <= 16'h0000;
      coeffs_in_data_log_force[1498] <= 16'h0000;
      coeffs_in_data_log_force[1499] <= 16'h0000;
      coeffs_in_data_log_force[1500] <= 16'h0000;
      coeffs_in_data_log_force[1501] <= 16'h0000;
      coeffs_in_data_log_force[1502] <= 16'h0000;
      coeffs_in_data_log_force[1503] <= 16'h0000;
      coeffs_in_data_log_force[1504] <= 16'h0000;
      coeffs_in_data_log_force[1505] <= 16'h0000;
      coeffs_in_data_log_force[1506] <= 16'h0000;
      coeffs_in_data_log_force[1507] <= 16'h0000;
      coeffs_in_data_log_force[1508] <= 16'h0000;
      coeffs_in_data_log_force[1509] <= 16'h0000;
      coeffs_in_data_log_force[1510] <= 16'h0000;
      coeffs_in_data_log_force[1511] <= 16'h0000;
      coeffs_in_data_log_force[1512] <= 16'h0000;
      coeffs_in_data_log_force[1513] <= 16'h0000;
      coeffs_in_data_log_force[1514] <= 16'h0000;
      coeffs_in_data_log_force[1515] <= 16'h0000;
      coeffs_in_data_log_force[1516] <= 16'h0000;
      coeffs_in_data_log_force[1517] <= 16'h0000;
      coeffs_in_data_log_force[1518] <= 16'h0000;
      coeffs_in_data_log_force[1519] <= 16'h0000;
      coeffs_in_data_log_force[1520] <= 16'h0000;
      coeffs_in_data_log_force[1521] <= 16'h0000;
      coeffs_in_data_log_force[1522] <= 16'h0000;
      coeffs_in_data_log_force[1523] <= 16'h0000;
      coeffs_in_data_log_force[1524] <= 16'h0000;
      coeffs_in_data_log_force[1525] <= 16'h0000;
      coeffs_in_data_log_force[1526] <= 16'h0000;
      coeffs_in_data_log_force[1527] <= 16'h0000;
      coeffs_in_data_log_force[1528] <= 16'h0000;
      coeffs_in_data_log_force[1529] <= 16'h0000;
      coeffs_in_data_log_force[1530] <= 16'h0000;
      coeffs_in_data_log_force[1531] <= 16'h0000;
      coeffs_in_data_log_force[1532] <= 16'h0000;
      coeffs_in_data_log_force[1533] <= 16'h0000;
      coeffs_in_data_log_force[1534] <= 16'h0000;
      coeffs_in_data_log_force[1535] <= 16'h0000;
      coeffs_in_data_log_force[1536] <= 16'h0000;
      coeffs_in_data_log_force[1537] <= 16'h0000;
      coeffs_in_data_log_force[1538] <= 16'h0000;
      coeffs_in_data_log_force[1539] <= 16'h0000;
      coeffs_in_data_log_force[1540] <= 16'h0000;
      coeffs_in_data_log_force[1541] <= 16'h0000;
      coeffs_in_data_log_force[1542] <= 16'h0000;
      coeffs_in_data_log_force[1543] <= 16'h0000;
      coeffs_in_data_log_force[1544] <= 16'h0000;
      coeffs_in_data_log_force[1545] <= 16'h0000;
      coeffs_in_data_log_force[1546] <= 16'h0000;
      coeffs_in_data_log_force[1547] <= 16'h0000;
      coeffs_in_data_log_force[1548] <= 16'h0000;
      coeffs_in_data_log_force[1549] <= 16'h0000;
      coeffs_in_data_log_force[1550] <= 16'h0000;
      coeffs_in_data_log_force[1551] <= 16'h0000;
      coeffs_in_data_log_force[1552] <= 16'h0000;
      coeffs_in_data_log_force[1553] <= 16'h0000;
      coeffs_in_data_log_force[1554] <= 16'h0000;
      coeffs_in_data_log_force[1555] <= 16'h0000;
      coeffs_in_data_log_force[1556] <= 16'h0000;
      coeffs_in_data_log_force[1557] <= 16'h0000;
      coeffs_in_data_log_force[1558] <= 16'h0000;
      coeffs_in_data_log_force[1559] <= 16'h0000;
      coeffs_in_data_log_force[1560] <= 16'h0000;
      coeffs_in_data_log_force[1561] <= 16'h0000;
      coeffs_in_data_log_force[1562] <= 16'h0000;
      coeffs_in_data_log_force[1563] <= 16'h0000;
      coeffs_in_data_log_force[1564] <= 16'h0000;
      coeffs_in_data_log_force[1565] <= 16'h0000;
      coeffs_in_data_log_force[1566] <= 16'h0000;
      coeffs_in_data_log_force[1567] <= 16'h0000;
      coeffs_in_data_log_force[1568] <= 16'h0000;
      coeffs_in_data_log_force[1569] <= 16'h0000;
      coeffs_in_data_log_force[1570] <= 16'h0000;
      coeffs_in_data_log_force[1571] <= 16'h0000;
      coeffs_in_data_log_force[1572] <= 16'h0000;
      coeffs_in_data_log_force[1573] <= 16'h0000;
      coeffs_in_data_log_force[1574] <= 16'h0000;
      coeffs_in_data_log_force[1575] <= 16'h0000;
      coeffs_in_data_log_force[1576] <= 16'h0000;
      coeffs_in_data_log_force[1577] <= 16'h0000;
      coeffs_in_data_log_force[1578] <= 16'h0000;
      coeffs_in_data_log_force[1579] <= 16'h0000;
      coeffs_in_data_log_force[1580] <= 16'h0000;
      coeffs_in_data_log_force[1581] <= 16'h0000;
      coeffs_in_data_log_force[1582] <= 16'h0000;
      coeffs_in_data_log_force[1583] <= 16'h0000;
      coeffs_in_data_log_force[1584] <= 16'h0000;
      coeffs_in_data_log_force[1585] <= 16'h0000;
      coeffs_in_data_log_force[1586] <= 16'h0000;
      coeffs_in_data_log_force[1587] <= 16'h0000;
      coeffs_in_data_log_force[1588] <= 16'h0000;
      coeffs_in_data_log_force[1589] <= 16'h0000;
      coeffs_in_data_log_force[1590] <= 16'h0000;
      coeffs_in_data_log_force[1591] <= 16'h0000;
      coeffs_in_data_log_force[1592] <= 16'h0000;
      coeffs_in_data_log_force[1593] <= 16'h0000;
      coeffs_in_data_log_force[1594] <= 16'h0000;
      coeffs_in_data_log_force[1595] <= 16'h0000;
      coeffs_in_data_log_force[1596] <= 16'h0000;
      coeffs_in_data_log_force[1597] <= 16'h0000;
      coeffs_in_data_log_force[1598] <= 16'h0000;
      coeffs_in_data_log_force[1599] <= 16'h0000;
      coeffs_in_data_log_force[1600] <= 16'h0000;
      coeffs_in_data_log_force[1601] <= 16'h0000;
      coeffs_in_data_log_force[1602] <= 16'h0000;
      coeffs_in_data_log_force[1603] <= 16'h0000;
      coeffs_in_data_log_force[1604] <= 16'h0000;
      coeffs_in_data_log_force[1605] <= 16'h0000;
      coeffs_in_data_log_force[1606] <= 16'h0000;
      coeffs_in_data_log_force[1607] <= 16'h0000;
      coeffs_in_data_log_force[1608] <= 16'h0000;
      coeffs_in_data_log_force[1609] <= 16'h0000;
      coeffs_in_data_log_force[1610] <= 16'h0000;
      coeffs_in_data_log_force[1611] <= 16'h0000;
      coeffs_in_data_log_force[1612] <= 16'h0000;
      coeffs_in_data_log_force[1613] <= 16'h0000;
      coeffs_in_data_log_force[1614] <= 16'h0000;
      coeffs_in_data_log_force[1615] <= 16'h0000;
      coeffs_in_data_log_force[1616] <= 16'h0000;
      coeffs_in_data_log_force[1617] <= 16'h0000;
      coeffs_in_data_log_force[1618] <= 16'h0000;
      coeffs_in_data_log_force[1619] <= 16'h0000;
      coeffs_in_data_log_force[1620] <= 16'h0000;
      coeffs_in_data_log_force[1621] <= 16'h0000;
      coeffs_in_data_log_force[1622] <= 16'h0000;
      coeffs_in_data_log_force[1623] <= 16'h0000;
      coeffs_in_data_log_force[1624] <= 16'h0000;
      coeffs_in_data_log_force[1625] <= 16'h0000;
      coeffs_in_data_log_force[1626] <= 16'h0000;
      coeffs_in_data_log_force[1627] <= 16'h0000;
      coeffs_in_data_log_force[1628] <= 16'h0000;
      coeffs_in_data_log_force[1629] <= 16'h0000;
      coeffs_in_data_log_force[1630] <= 16'h0000;
      coeffs_in_data_log_force[1631] <= 16'h0000;
      coeffs_in_data_log_force[1632] <= 16'h0000;
      coeffs_in_data_log_force[1633] <= 16'h0000;
      coeffs_in_data_log_force[1634] <= 16'h0000;
      coeffs_in_data_log_force[1635] <= 16'h0000;
      coeffs_in_data_log_force[1636] <= 16'h0000;
      coeffs_in_data_log_force[1637] <= 16'h0000;
      coeffs_in_data_log_force[1638] <= 16'h0000;
      coeffs_in_data_log_force[1639] <= 16'h0000;
      coeffs_in_data_log_force[1640] <= 16'h0000;
      coeffs_in_data_log_force[1641] <= 16'h0000;
      coeffs_in_data_log_force[1642] <= 16'h0000;
      coeffs_in_data_log_force[1643] <= 16'h0000;
      coeffs_in_data_log_force[1644] <= 16'h0000;
      coeffs_in_data_log_force[1645] <= 16'h0000;
      coeffs_in_data_log_force[1646] <= 16'h0000;
      coeffs_in_data_log_force[1647] <= 16'h0000;
      coeffs_in_data_log_force[1648] <= 16'h0000;
      coeffs_in_data_log_force[1649] <= 16'h0000;
      coeffs_in_data_log_force[1650] <= 16'h0000;
      coeffs_in_data_log_force[1651] <= 16'h0000;
      coeffs_in_data_log_force[1652] <= 16'h0000;
      coeffs_in_data_log_force[1653] <= 16'h0000;
      coeffs_in_data_log_force[1654] <= 16'h0000;
      coeffs_in_data_log_force[1655] <= 16'h0000;
      coeffs_in_data_log_force[1656] <= 16'h0000;
      coeffs_in_data_log_force[1657] <= 16'h0000;
      coeffs_in_data_log_force[1658] <= 16'h0000;
      coeffs_in_data_log_force[1659] <= 16'h0000;
      coeffs_in_data_log_force[1660] <= 16'h0000;
      coeffs_in_data_log_force[1661] <= 16'h0000;
      coeffs_in_data_log_force[1662] <= 16'h0000;
      coeffs_in_data_log_force[1663] <= 16'h0000;
      coeffs_in_data_log_force[1664] <= 16'h0000;
      coeffs_in_data_log_force[1665] <= 16'h0000;
      coeffs_in_data_log_force[1666] <= 16'h0000;
      coeffs_in_data_log_force[1667] <= 16'h0000;
      coeffs_in_data_log_force[1668] <= 16'h0000;
      coeffs_in_data_log_force[1669] <= 16'h0000;
      coeffs_in_data_log_force[1670] <= 16'h0000;
      coeffs_in_data_log_force[1671] <= 16'h0000;
      coeffs_in_data_log_force[1672] <= 16'h0000;
      coeffs_in_data_log_force[1673] <= 16'h0000;
      coeffs_in_data_log_force[1674] <= 16'h0000;
      coeffs_in_data_log_force[1675] <= 16'h0000;
      coeffs_in_data_log_force[1676] <= 16'h0000;
      coeffs_in_data_log_force[1677] <= 16'h0000;
      coeffs_in_data_log_force[1678] <= 16'h0000;
      coeffs_in_data_log_force[1679] <= 16'h0000;
      coeffs_in_data_log_force[1680] <= 16'h0000;
      coeffs_in_data_log_force[1681] <= 16'h0000;
      coeffs_in_data_log_force[1682] <= 16'h0000;
      coeffs_in_data_log_force[1683] <= 16'h0000;
      coeffs_in_data_log_force[1684] <= 16'h0000;
      coeffs_in_data_log_force[1685] <= 16'h0000;
      coeffs_in_data_log_force[1686] <= 16'h0000;
      coeffs_in_data_log_force[1687] <= 16'h0000;
      coeffs_in_data_log_force[1688] <= 16'h0000;
      coeffs_in_data_log_force[1689] <= 16'h0000;
      coeffs_in_data_log_force[1690] <= 16'h0000;
      coeffs_in_data_log_force[1691] <= 16'h0000;
      coeffs_in_data_log_force[1692] <= 16'h0000;
      coeffs_in_data_log_force[1693] <= 16'h0000;
      coeffs_in_data_log_force[1694] <= 16'h0000;
      coeffs_in_data_log_force[1695] <= 16'h0000;
      coeffs_in_data_log_force[1696] <= 16'h0000;
      coeffs_in_data_log_force[1697] <= 16'h0000;
      coeffs_in_data_log_force[1698] <= 16'h0000;
      coeffs_in_data_log_force[1699] <= 16'h0000;
      coeffs_in_data_log_force[1700] <= 16'h0000;
      coeffs_in_data_log_force[1701] <= 16'h0000;
      coeffs_in_data_log_force[1702] <= 16'h0000;
      coeffs_in_data_log_force[1703] <= 16'h0000;
      coeffs_in_data_log_force[1704] <= 16'h0000;
      coeffs_in_data_log_force[1705] <= 16'h0000;
      coeffs_in_data_log_force[1706] <= 16'h0000;
      coeffs_in_data_log_force[1707] <= 16'h0000;
      coeffs_in_data_log_force[1708] <= 16'h0000;
      coeffs_in_data_log_force[1709] <= 16'h0000;
      coeffs_in_data_log_force[1710] <= 16'h0000;
      coeffs_in_data_log_force[1711] <= 16'h0000;
      coeffs_in_data_log_force[1712] <= 16'h0000;
      coeffs_in_data_log_force[1713] <= 16'h0000;
      coeffs_in_data_log_force[1714] <= 16'h0000;
      coeffs_in_data_log_force[1715] <= 16'h0000;
      coeffs_in_data_log_force[1716] <= 16'h0000;
      coeffs_in_data_log_force[1717] <= 16'h0000;
      coeffs_in_data_log_force[1718] <= 16'h0000;
      coeffs_in_data_log_force[1719] <= 16'h0000;
      coeffs_in_data_log_force[1720] <= 16'h0000;
      coeffs_in_data_log_force[1721] <= 16'h0000;
      coeffs_in_data_log_force[1722] <= 16'h0000;
      coeffs_in_data_log_force[1723] <= 16'h0000;
      coeffs_in_data_log_force[1724] <= 16'h0000;
      coeffs_in_data_log_force[1725] <= 16'h0000;
      coeffs_in_data_log_force[1726] <= 16'h0000;
      coeffs_in_data_log_force[1727] <= 16'h0000;
      coeffs_in_data_log_force[1728] <= 16'h0000;
      coeffs_in_data_log_force[1729] <= 16'h0000;
      coeffs_in_data_log_force[1730] <= 16'h0000;
      coeffs_in_data_log_force[1731] <= 16'h0000;
      coeffs_in_data_log_force[1732] <= 16'h0000;
      coeffs_in_data_log_force[1733] <= 16'h0000;
      coeffs_in_data_log_force[1734] <= 16'h0000;
      coeffs_in_data_log_force[1735] <= 16'h0000;
      coeffs_in_data_log_force[1736] <= 16'h0000;
      coeffs_in_data_log_force[1737] <= 16'h0000;
      coeffs_in_data_log_force[1738] <= 16'h0000;
      coeffs_in_data_log_force[1739] <= 16'h0000;
      coeffs_in_data_log_force[1740] <= 16'h0000;
      coeffs_in_data_log_force[1741] <= 16'h0000;
      coeffs_in_data_log_force[1742] <= 16'h0000;
      coeffs_in_data_log_force[1743] <= 16'h0000;
      coeffs_in_data_log_force[1744] <= 16'h0000;
      coeffs_in_data_log_force[1745] <= 16'h0000;
      coeffs_in_data_log_force[1746] <= 16'h0000;
      coeffs_in_data_log_force[1747] <= 16'h0000;
      coeffs_in_data_log_force[1748] <= 16'h0000;
      coeffs_in_data_log_force[1749] <= 16'h0000;
      coeffs_in_data_log_force[1750] <= 16'h0000;
      coeffs_in_data_log_force[1751] <= 16'h0000;
      coeffs_in_data_log_force[1752] <= 16'h0000;
      coeffs_in_data_log_force[1753] <= 16'h0000;
      coeffs_in_data_log_force[1754] <= 16'h0000;
      coeffs_in_data_log_force[1755] <= 16'h0000;
      coeffs_in_data_log_force[1756] <= 16'h0000;
      coeffs_in_data_log_force[1757] <= 16'h0000;
      coeffs_in_data_log_force[1758] <= 16'h0000;
      coeffs_in_data_log_force[1759] <= 16'h0000;
      coeffs_in_data_log_force[1760] <= 16'h0000;
      coeffs_in_data_log_force[1761] <= 16'h0000;
      coeffs_in_data_log_force[1762] <= 16'h0000;
      coeffs_in_data_log_force[1763] <= 16'h0000;
      coeffs_in_data_log_force[1764] <= 16'h0000;
      coeffs_in_data_log_force[1765] <= 16'h0000;
      coeffs_in_data_log_force[1766] <= 16'h0000;
      coeffs_in_data_log_force[1767] <= 16'h0000;
      coeffs_in_data_log_force[1768] <= 16'h0000;
      coeffs_in_data_log_force[1769] <= 16'h0000;
      coeffs_in_data_log_force[1770] <= 16'h0000;
      coeffs_in_data_log_force[1771] <= 16'h0000;
      coeffs_in_data_log_force[1772] <= 16'h0000;
      coeffs_in_data_log_force[1773] <= 16'h0000;
      coeffs_in_data_log_force[1774] <= 16'h0000;
      coeffs_in_data_log_force[1775] <= 16'h0000;
      coeffs_in_data_log_force[1776] <= 16'h0000;
      coeffs_in_data_log_force[1777] <= 16'h0000;
      coeffs_in_data_log_force[1778] <= 16'h0000;
      coeffs_in_data_log_force[1779] <= 16'h0000;
      coeffs_in_data_log_force[1780] <= 16'h0000;
      coeffs_in_data_log_force[1781] <= 16'h0000;
      coeffs_in_data_log_force[1782] <= 16'h0000;
      coeffs_in_data_log_force[1783] <= 16'h0000;
      coeffs_in_data_log_force[1784] <= 16'h0000;
      coeffs_in_data_log_force[1785] <= 16'h0000;
      coeffs_in_data_log_force[1786] <= 16'h0000;
      coeffs_in_data_log_force[1787] <= 16'h0000;
      coeffs_in_data_log_force[1788] <= 16'h0000;
      coeffs_in_data_log_force[1789] <= 16'h0000;
      coeffs_in_data_log_force[1790] <= 16'h0000;
      coeffs_in_data_log_force[1791] <= 16'h0000;
      coeffs_in_data_log_force[1792] <= 16'h0000;
      coeffs_in_data_log_force[1793] <= 16'h0000;
      coeffs_in_data_log_force[1794] <= 16'h0000;
      coeffs_in_data_log_force[1795] <= 16'h0000;
      coeffs_in_data_log_force[1796] <= 16'h0000;
      coeffs_in_data_log_force[1797] <= 16'h0000;
      coeffs_in_data_log_force[1798] <= 16'h0000;
      coeffs_in_data_log_force[1799] <= 16'h0000;
      coeffs_in_data_log_force[1800] <= 16'h0000;
      coeffs_in_data_log_force[1801] <= 16'h0000;
      coeffs_in_data_log_force[1802] <= 16'h0000;
      coeffs_in_data_log_force[1803] <= 16'h0000;
      coeffs_in_data_log_force[1804] <= 16'h0000;
      coeffs_in_data_log_force[1805] <= 16'h0000;
      coeffs_in_data_log_force[1806] <= 16'h0000;
      coeffs_in_data_log_force[1807] <= 16'h0000;
      coeffs_in_data_log_force[1808] <= 16'h0000;
      coeffs_in_data_log_force[1809] <= 16'h0000;
      coeffs_in_data_log_force[1810] <= 16'h0000;
      coeffs_in_data_log_force[1811] <= 16'h0000;
      coeffs_in_data_log_force[1812] <= 16'h0000;
      coeffs_in_data_log_force[1813] <= 16'h0000;
      coeffs_in_data_log_force[1814] <= 16'h0000;
      coeffs_in_data_log_force[1815] <= 16'h0000;
      coeffs_in_data_log_force[1816] <= 16'h0000;
      coeffs_in_data_log_force[1817] <= 16'h0000;
      coeffs_in_data_log_force[1818] <= 16'h0000;
      coeffs_in_data_log_force[1819] <= 16'h0000;
      coeffs_in_data_log_force[1820] <= 16'h0000;
      coeffs_in_data_log_force[1821] <= 16'h0000;
      coeffs_in_data_log_force[1822] <= 16'h0000;
      coeffs_in_data_log_force[1823] <= 16'h0000;
      coeffs_in_data_log_force[1824] <= 16'h0000;
      coeffs_in_data_log_force[1825] <= 16'h0000;
      coeffs_in_data_log_force[1826] <= 16'h0000;
      coeffs_in_data_log_force[1827] <= 16'h0000;
      coeffs_in_data_log_force[1828] <= 16'h0000;
      coeffs_in_data_log_force[1829] <= 16'h0000;
      coeffs_in_data_log_force[1830] <= 16'h0000;
      coeffs_in_data_log_force[1831] <= 16'h0000;
      coeffs_in_data_log_force[1832] <= 16'h0000;
      coeffs_in_data_log_force[1833] <= 16'h0000;
      coeffs_in_data_log_force[1834] <= 16'h0000;
      coeffs_in_data_log_force[1835] <= 16'h0000;
      coeffs_in_data_log_force[1836] <= 16'h0000;
      coeffs_in_data_log_force[1837] <= 16'h0000;
      coeffs_in_data_log_force[1838] <= 16'h0000;
      coeffs_in_data_log_force[1839] <= 16'h0000;
      coeffs_in_data_log_force[1840] <= 16'h0000;
      coeffs_in_data_log_force[1841] <= 16'h0000;
      coeffs_in_data_log_force[1842] <= 16'h0000;
      coeffs_in_data_log_force[1843] <= 16'h0000;
      coeffs_in_data_log_force[1844] <= 16'h0000;
      coeffs_in_data_log_force[1845] <= 16'h0000;
      coeffs_in_data_log_force[1846] <= 16'h0000;
      coeffs_in_data_log_force[1847] <= 16'h0000;
      coeffs_in_data_log_force[1848] <= 16'h0000;
      coeffs_in_data_log_force[1849] <= 16'h0000;
      coeffs_in_data_log_force[1850] <= 16'h0000;
      coeffs_in_data_log_force[1851] <= 16'h0000;
      coeffs_in_data_log_force[1852] <= 16'h0000;
      coeffs_in_data_log_force[1853] <= 16'h0000;
      coeffs_in_data_log_force[1854] <= 16'h0000;
      coeffs_in_data_log_force[1855] <= 16'h0000;
      coeffs_in_data_log_force[1856] <= 16'h0000;
      coeffs_in_data_log_force[1857] <= 16'h0000;
      coeffs_in_data_log_force[1858] <= 16'h0000;
      coeffs_in_data_log_force[1859] <= 16'h0000;
      coeffs_in_data_log_force[1860] <= 16'h0000;
      coeffs_in_data_log_force[1861] <= 16'h0000;
      coeffs_in_data_log_force[1862] <= 16'h0000;
      coeffs_in_data_log_force[1863] <= 16'h0000;
      coeffs_in_data_log_force[1864] <= 16'h0000;
      coeffs_in_data_log_force[1865] <= 16'h0000;
      coeffs_in_data_log_force[1866] <= 16'h0000;
      coeffs_in_data_log_force[1867] <= 16'h0000;
      coeffs_in_data_log_force[1868] <= 16'h0000;
      coeffs_in_data_log_force[1869] <= 16'h0000;
      coeffs_in_data_log_force[1870] <= 16'h0000;
      coeffs_in_data_log_force[1871] <= 16'h0000;
      coeffs_in_data_log_force[1872] <= 16'h0000;
      coeffs_in_data_log_force[1873] <= 16'h0000;
      coeffs_in_data_log_force[1874] <= 16'h0000;
      coeffs_in_data_log_force[1875] <= 16'h0000;
      coeffs_in_data_log_force[1876] <= 16'h0000;
      coeffs_in_data_log_force[1877] <= 16'h0000;
      coeffs_in_data_log_force[1878] <= 16'h0000;
      coeffs_in_data_log_force[1879] <= 16'h0000;
      coeffs_in_data_log_force[1880] <= 16'h0000;
      coeffs_in_data_log_force[1881] <= 16'h0000;
      coeffs_in_data_log_force[1882] <= 16'h0000;
      coeffs_in_data_log_force[1883] <= 16'h0000;
      coeffs_in_data_log_force[1884] <= 16'h0000;
      coeffs_in_data_log_force[1885] <= 16'h0000;
      coeffs_in_data_log_force[1886] <= 16'h0000;
      coeffs_in_data_log_force[1887] <= 16'h0000;
      coeffs_in_data_log_force[1888] <= 16'h0000;
      coeffs_in_data_log_force[1889] <= 16'h0000;
      coeffs_in_data_log_force[1890] <= 16'h0000;
      coeffs_in_data_log_force[1891] <= 16'h0000;
      coeffs_in_data_log_force[1892] <= 16'h0000;
      coeffs_in_data_log_force[1893] <= 16'h0000;
      coeffs_in_data_log_force[1894] <= 16'h0000;
      coeffs_in_data_log_force[1895] <= 16'h0000;
      coeffs_in_data_log_force[1896] <= 16'h0000;
      coeffs_in_data_log_force[1897] <= 16'h0000;
      coeffs_in_data_log_force[1898] <= 16'h0000;
      coeffs_in_data_log_force[1899] <= 16'h0000;
      coeffs_in_data_log_force[1900] <= 16'h0000;
      coeffs_in_data_log_force[1901] <= 16'h0000;
      coeffs_in_data_log_force[1902] <= 16'h0000;
      coeffs_in_data_log_force[1903] <= 16'h0000;
      coeffs_in_data_log_force[1904] <= 16'h0000;
      coeffs_in_data_log_force[1905] <= 16'h0000;
      coeffs_in_data_log_force[1906] <= 16'h0000;
      coeffs_in_data_log_force[1907] <= 16'h0000;
      coeffs_in_data_log_force[1908] <= 16'h0000;
      coeffs_in_data_log_force[1909] <= 16'h0000;
      coeffs_in_data_log_force[1910] <= 16'h0000;
      coeffs_in_data_log_force[1911] <= 16'h0000;
      coeffs_in_data_log_force[1912] <= 16'h0000;
      coeffs_in_data_log_force[1913] <= 16'h0000;
      coeffs_in_data_log_force[1914] <= 16'h0000;
      coeffs_in_data_log_force[1915] <= 16'h0000;
      coeffs_in_data_log_force[1916] <= 16'h0000;
      coeffs_in_data_log_force[1917] <= 16'h0000;
      coeffs_in_data_log_force[1918] <= 16'h0000;
      coeffs_in_data_log_force[1919] <= 16'h0000;
      coeffs_in_data_log_force[1920] <= 16'h0000;
      coeffs_in_data_log_force[1921] <= 16'h0000;
      coeffs_in_data_log_force[1922] <= 16'h0000;
      coeffs_in_data_log_force[1923] <= 16'h0000;
      coeffs_in_data_log_force[1924] <= 16'h0000;
      coeffs_in_data_log_force[1925] <= 16'h0000;
      coeffs_in_data_log_force[1926] <= 16'h0000;
      coeffs_in_data_log_force[1927] <= 16'h0000;
      coeffs_in_data_log_force[1928] <= 16'h0000;
      coeffs_in_data_log_force[1929] <= 16'h0000;
      coeffs_in_data_log_force[1930] <= 16'h0000;
      coeffs_in_data_log_force[1931] <= 16'h0000;
      coeffs_in_data_log_force[1932] <= 16'h0000;
      coeffs_in_data_log_force[1933] <= 16'h0000;
      coeffs_in_data_log_force[1934] <= 16'h0000;
      coeffs_in_data_log_force[1935] <= 16'h0000;
      coeffs_in_data_log_force[1936] <= 16'h0000;
      coeffs_in_data_log_force[1937] <= 16'h0000;
      coeffs_in_data_log_force[1938] <= 16'h0000;
      coeffs_in_data_log_force[1939] <= 16'h0000;
      coeffs_in_data_log_force[1940] <= 16'h0000;
      coeffs_in_data_log_force[1941] <= 16'h0000;
      coeffs_in_data_log_force[1942] <= 16'h0000;
      coeffs_in_data_log_force[1943] <= 16'h0000;
      coeffs_in_data_log_force[1944] <= 16'h0000;
      coeffs_in_data_log_force[1945] <= 16'h0000;
      coeffs_in_data_log_force[1946] <= 16'h0000;
      coeffs_in_data_log_force[1947] <= 16'h0000;
      coeffs_in_data_log_force[1948] <= 16'h0000;
      coeffs_in_data_log_force[1949] <= 16'h0000;
      coeffs_in_data_log_force[1950] <= 16'h0000;
      coeffs_in_data_log_force[1951] <= 16'h0000;
      coeffs_in_data_log_force[1952] <= 16'h0000;
      coeffs_in_data_log_force[1953] <= 16'h0000;
      coeffs_in_data_log_force[1954] <= 16'h0000;
      coeffs_in_data_log_force[1955] <= 16'h0000;
      coeffs_in_data_log_force[1956] <= 16'h0000;
      coeffs_in_data_log_force[1957] <= 16'h0000;
      coeffs_in_data_log_force[1958] <= 16'h0000;
      coeffs_in_data_log_force[1959] <= 16'h0000;
      coeffs_in_data_log_force[1960] <= 16'h0000;
      coeffs_in_data_log_force[1961] <= 16'h0000;
      coeffs_in_data_log_force[1962] <= 16'h0000;
      coeffs_in_data_log_force[1963] <= 16'h0000;
      coeffs_in_data_log_force[1964] <= 16'h0000;
      coeffs_in_data_log_force[1965] <= 16'h0000;
      coeffs_in_data_log_force[1966] <= 16'h0000;
      coeffs_in_data_log_force[1967] <= 16'h0000;
      coeffs_in_data_log_force[1968] <= 16'h0000;
      coeffs_in_data_log_force[1969] <= 16'h0000;
      coeffs_in_data_log_force[1970] <= 16'h0000;
      coeffs_in_data_log_force[1971] <= 16'h0000;
      coeffs_in_data_log_force[1972] <= 16'h0000;
      coeffs_in_data_log_force[1973] <= 16'h0000;
      coeffs_in_data_log_force[1974] <= 16'h0000;
      coeffs_in_data_log_force[1975] <= 16'h0000;
      coeffs_in_data_log_force[1976] <= 16'h0000;
      coeffs_in_data_log_force[1977] <= 16'h0000;
      coeffs_in_data_log_force[1978] <= 16'h0000;
      coeffs_in_data_log_force[1979] <= 16'h0000;
      coeffs_in_data_log_force[1980] <= 16'h0000;
      coeffs_in_data_log_force[1981] <= 16'h0000;
      coeffs_in_data_log_force[1982] <= 16'h0000;
      coeffs_in_data_log_force[1983] <= 16'h0000;
      coeffs_in_data_log_force[1984] <= 16'h0000;
      coeffs_in_data_log_force[1985] <= 16'h0000;
      coeffs_in_data_log_force[1986] <= 16'h0000;
      coeffs_in_data_log_force[1987] <= 16'h0000;
      coeffs_in_data_log_force[1988] <= 16'h0000;
      coeffs_in_data_log_force[1989] <= 16'h0000;
      coeffs_in_data_log_force[1990] <= 16'h0000;
      coeffs_in_data_log_force[1991] <= 16'h0000;
      coeffs_in_data_log_force[1992] <= 16'h0000;
      coeffs_in_data_log_force[1993] <= 16'h0000;
      coeffs_in_data_log_force[1994] <= 16'h0000;
      coeffs_in_data_log_force[1995] <= 16'h0000;
      coeffs_in_data_log_force[1996] <= 16'h0000;
      coeffs_in_data_log_force[1997] <= 16'h0000;
      coeffs_in_data_log_force[1998] <= 16'h0000;
      coeffs_in_data_log_force[1999] <= 16'h0000;
      coeffs_in_data_log_force[2000] <= 16'h0000;
      coeffs_in_data_log_force[2001] <= 16'h0000;
      coeffs_in_data_log_force[2002] <= 16'h0000;
      coeffs_in_data_log_force[2003] <= 16'h0000;
      coeffs_in_data_log_force[2004] <= 16'h0000;
      coeffs_in_data_log_force[2005] <= 16'h0000;
      coeffs_in_data_log_force[2006] <= 16'h0000;
      coeffs_in_data_log_force[2007] <= 16'h0000;
      coeffs_in_data_log_force[2008] <= 16'h0000;
      coeffs_in_data_log_force[2009] <= 16'h0000;
      coeffs_in_data_log_force[2010] <= 16'h0000;
      coeffs_in_data_log_force[2011] <= 16'h0000;
      coeffs_in_data_log_force[2012] <= 16'h0000;
      coeffs_in_data_log_force[2013] <= 16'h0000;
      coeffs_in_data_log_force[2014] <= 16'h0000;
      coeffs_in_data_log_force[2015] <= 16'h0000;
      coeffs_in_data_log_force[2016] <= 16'h0000;
      coeffs_in_data_log_force[2017] <= 16'h0000;
      coeffs_in_data_log_force[2018] <= 16'h0000;
      coeffs_in_data_log_force[2019] <= 16'h0000;
      coeffs_in_data_log_force[2020] <= 16'h0000;
      coeffs_in_data_log_force[2021] <= 16'h0000;
      coeffs_in_data_log_force[2022] <= 16'h0000;
      coeffs_in_data_log_force[2023] <= 16'h0000;
      coeffs_in_data_log_force[2024] <= 16'h0000;
      coeffs_in_data_log_force[2025] <= 16'h0000;
      coeffs_in_data_log_force[2026] <= 16'h0000;
      coeffs_in_data_log_force[2027] <= 16'h0000;
      coeffs_in_data_log_force[2028] <= 16'h0000;
      coeffs_in_data_log_force[2029] <= 16'h0000;
      coeffs_in_data_log_force[2030] <= 16'h0000;
      coeffs_in_data_log_force[2031] <= 16'h0000;
      coeffs_in_data_log_force[2032] <= 16'h0000;
      coeffs_in_data_log_force[2033] <= 16'h0000;
      coeffs_in_data_log_force[2034] <= 16'h0000;
      coeffs_in_data_log_force[2035] <= 16'h0000;
      coeffs_in_data_log_force[2036] <= 16'h0000;
      coeffs_in_data_log_force[2037] <= 16'h0000;
      coeffs_in_data_log_force[2038] <= 16'h0000;
      coeffs_in_data_log_force[2039] <= 16'h0000;
      coeffs_in_data_log_force[2040] <= 16'h0000;
      coeffs_in_data_log_force[2041] <= 16'h0000;
      coeffs_in_data_log_force[2042] <= 16'h0000;
      coeffs_in_data_log_force[2043] <= 16'h0000;
      coeffs_in_data_log_force[2044] <= 16'h0000;
      coeffs_in_data_log_force[2045] <= 16'h0000;
      coeffs_in_data_log_force[2046] <= 16'h0000;
      coeffs_in_data_log_force[2047] <= 16'h0000;
      coeffs_in_data_log_force[2048] <= 16'h0000;
      coeffs_in_data_log_force[2049] <= 16'h0000;
      coeffs_in_data_log_force[2050] <= 16'h0000;
      coeffs_in_data_log_force[2051] <= 16'h0000;
      coeffs_in_data_log_force[2052] <= 16'h0000;
      coeffs_in_data_log_force[2053] <= 16'h0000;
      coeffs_in_data_log_force[2054] <= 16'h0000;
      coeffs_in_data_log_force[2055] <= 16'h0000;
      coeffs_in_data_log_force[2056] <= 16'h0000;
      coeffs_in_data_log_force[2057] <= 16'h0000;
      coeffs_in_data_log_force[2058] <= 16'h0000;
      coeffs_in_data_log_force[2059] <= 16'h0000;
      coeffs_in_data_log_force[2060] <= 16'h0000;
      coeffs_in_data_log_force[2061] <= 16'h0000;
      coeffs_in_data_log_force[2062] <= 16'h0000;
      coeffs_in_data_log_force[2063] <= 16'h0000;
      coeffs_in_data_log_force[2064] <= 16'h0000;
      coeffs_in_data_log_force[2065] <= 16'h0000;
      coeffs_in_data_log_force[2066] <= 16'h0000;
      coeffs_in_data_log_force[2067] <= 16'h0000;
      coeffs_in_data_log_force[2068] <= 16'h0000;
      coeffs_in_data_log_force[2069] <= 16'h0000;
      coeffs_in_data_log_force[2070] <= 16'h0000;
      coeffs_in_data_log_force[2071] <= 16'h0000;
      coeffs_in_data_log_force[2072] <= 16'h0000;
      coeffs_in_data_log_force[2073] <= 16'h0000;
      coeffs_in_data_log_force[2074] <= 16'h0000;
      coeffs_in_data_log_force[2075] <= 16'h0000;
      coeffs_in_data_log_force[2076] <= 16'h0000;
      coeffs_in_data_log_force[2077] <= 16'h0000;
      coeffs_in_data_log_force[2078] <= 16'h0000;
      coeffs_in_data_log_force[2079] <= 16'h0000;
      coeffs_in_data_log_force[2080] <= 16'h0000;
      coeffs_in_data_log_force[2081] <= 16'h0000;
      coeffs_in_data_log_force[2082] <= 16'h0000;
      coeffs_in_data_log_force[2083] <= 16'h0000;
      coeffs_in_data_log_force[2084] <= 16'h0000;
      coeffs_in_data_log_force[2085] <= 16'h0000;
      coeffs_in_data_log_force[2086] <= 16'h0000;
      coeffs_in_data_log_force[2087] <= 16'h0000;
      coeffs_in_data_log_force[2088] <= 16'h0000;
      coeffs_in_data_log_force[2089] <= 16'h0000;
      coeffs_in_data_log_force[2090] <= 16'h0000;
      coeffs_in_data_log_force[2091] <= 16'h0000;
      coeffs_in_data_log_force[2092] <= 16'h0000;
      coeffs_in_data_log_force[2093] <= 16'h0000;
      coeffs_in_data_log_force[2094] <= 16'h0000;
      coeffs_in_data_log_force[2095] <= 16'h0000;
      coeffs_in_data_log_force[2096] <= 16'h0000;
      coeffs_in_data_log_force[2097] <= 16'h0000;
      coeffs_in_data_log_force[2098] <= 16'h0000;
      coeffs_in_data_log_force[2099] <= 16'h0000;
      coeffs_in_data_log_force[2100] <= 16'h0000;
      coeffs_in_data_log_force[2101] <= 16'h0000;
      coeffs_in_data_log_force[2102] <= 16'h0000;
      coeffs_in_data_log_force[2103] <= 16'h0000;
      coeffs_in_data_log_force[2104] <= 16'h0000;
      coeffs_in_data_log_force[2105] <= 16'h0000;
      coeffs_in_data_log_force[2106] <= 16'h0000;
      coeffs_in_data_log_force[2107] <= 16'h0000;
      coeffs_in_data_log_force[2108] <= 16'h0000;
      coeffs_in_data_log_force[2109] <= 16'h0000;
      coeffs_in_data_log_force[2110] <= 16'h0000;
      coeffs_in_data_log_force[2111] <= 16'h0000;
      coeffs_in_data_log_force[2112] <= 16'h0000;
      coeffs_in_data_log_force[2113] <= 16'h0000;
      coeffs_in_data_log_force[2114] <= 16'h0000;
      coeffs_in_data_log_force[2115] <= 16'h0000;
      coeffs_in_data_log_force[2116] <= 16'h0000;
      coeffs_in_data_log_force[2117] <= 16'h0000;
      coeffs_in_data_log_force[2118] <= 16'h0000;
      coeffs_in_data_log_force[2119] <= 16'h0000;
      coeffs_in_data_log_force[2120] <= 16'h0000;
      coeffs_in_data_log_force[2121] <= 16'h0000;
      coeffs_in_data_log_force[2122] <= 16'h0000;
      coeffs_in_data_log_force[2123] <= 16'h0000;
      coeffs_in_data_log_force[2124] <= 16'h0000;
      coeffs_in_data_log_force[2125] <= 16'h0000;
      coeffs_in_data_log_force[2126] <= 16'h0000;
      coeffs_in_data_log_force[2127] <= 16'h0000;
      coeffs_in_data_log_force[2128] <= 16'h0000;
      coeffs_in_data_log_force[2129] <= 16'h0000;
      coeffs_in_data_log_force[2130] <= 16'h0000;
      coeffs_in_data_log_force[2131] <= 16'h0000;
      coeffs_in_data_log_force[2132] <= 16'h0000;
      coeffs_in_data_log_force[2133] <= 16'h0000;
      coeffs_in_data_log_force[2134] <= 16'h0000;
      coeffs_in_data_log_force[2135] <= 16'h0000;
      coeffs_in_data_log_force[2136] <= 16'h0000;
      coeffs_in_data_log_force[2137] <= 16'h0000;
      coeffs_in_data_log_force[2138] <= 16'h0000;
      coeffs_in_data_log_force[2139] <= 16'h0000;
      coeffs_in_data_log_force[2140] <= 16'h0000;
      coeffs_in_data_log_force[2141] <= 16'h0000;
      coeffs_in_data_log_force[2142] <= 16'h0000;
      coeffs_in_data_log_force[2143] <= 16'h0000;
      coeffs_in_data_log_force[2144] <= 16'h0000;
      coeffs_in_data_log_force[2145] <= 16'h0000;
      coeffs_in_data_log_force[2146] <= 16'h0000;
      coeffs_in_data_log_force[2147] <= 16'h0000;
      coeffs_in_data_log_force[2148] <= 16'h0000;
      coeffs_in_data_log_force[2149] <= 16'h0000;
      coeffs_in_data_log_force[2150] <= 16'h0000;
      coeffs_in_data_log_force[2151] <= 16'h0000;
      coeffs_in_data_log_force[2152] <= 16'h0000;
      coeffs_in_data_log_force[2153] <= 16'h0000;
      coeffs_in_data_log_force[2154] <= 16'h0000;
      coeffs_in_data_log_force[2155] <= 16'h0000;
      coeffs_in_data_log_force[2156] <= 16'h0000;
      coeffs_in_data_log_force[2157] <= 16'h0000;
      coeffs_in_data_log_force[2158] <= 16'h0000;
      coeffs_in_data_log_force[2159] <= 16'h0000;
      coeffs_in_data_log_force[2160] <= 16'h0000;
      coeffs_in_data_log_force[2161] <= 16'h0000;
      coeffs_in_data_log_force[2162] <= 16'h0000;
      coeffs_in_data_log_force[2163] <= 16'h0000;
      coeffs_in_data_log_force[2164] <= 16'h0000;
      coeffs_in_data_log_force[2165] <= 16'h0000;
      coeffs_in_data_log_force[2166] <= 16'h0000;
      coeffs_in_data_log_force[2167] <= 16'h0000;
      coeffs_in_data_log_force[2168] <= 16'h0000;
      coeffs_in_data_log_force[2169] <= 16'h0000;
      coeffs_in_data_log_force[2170] <= 16'h0000;
      coeffs_in_data_log_force[2171] <= 16'h0000;
      coeffs_in_data_log_force[2172] <= 16'h0000;
      coeffs_in_data_log_force[2173] <= 16'h0000;
      coeffs_in_data_log_force[2174] <= 16'h0000;
      coeffs_in_data_log_force[2175] <= 16'h0000;
      coeffs_in_data_log_force[2176] <= 16'h0000;
      coeffs_in_data_log_force[2177] <= 16'h0000;
      coeffs_in_data_log_force[2178] <= 16'h0000;
      coeffs_in_data_log_force[2179] <= 16'h0000;
      coeffs_in_data_log_force[2180] <= 16'h0000;
      coeffs_in_data_log_force[2181] <= 16'h0000;
      coeffs_in_data_log_force[2182] <= 16'h0000;
      coeffs_in_data_log_force[2183] <= 16'h0000;
      coeffs_in_data_log_force[2184] <= 16'h0000;
      coeffs_in_data_log_force[2185] <= 16'h0000;
      coeffs_in_data_log_force[2186] <= 16'h0000;
      coeffs_in_data_log_force[2187] <= 16'h0000;
      coeffs_in_data_log_force[2188] <= 16'h0000;
      coeffs_in_data_log_force[2189] <= 16'h0000;
      coeffs_in_data_log_force[2190] <= 16'h0000;
      coeffs_in_data_log_force[2191] <= 16'h0000;
      coeffs_in_data_log_force[2192] <= 16'h0000;
      coeffs_in_data_log_force[2193] <= 16'h0000;
      coeffs_in_data_log_force[2194] <= 16'h0000;
      coeffs_in_data_log_force[2195] <= 16'h0000;
      coeffs_in_data_log_force[2196] <= 16'h0000;
      coeffs_in_data_log_force[2197] <= 16'h0000;
      coeffs_in_data_log_force[2198] <= 16'h0000;
      coeffs_in_data_log_force[2199] <= 16'h0000;
      coeffs_in_data_log_force[2200] <= 16'h0000;
      coeffs_in_data_log_force[2201] <= 16'h0000;
      coeffs_in_data_log_force[2202] <= 16'h0000;
      coeffs_in_data_log_force[2203] <= 16'h0000;
      coeffs_in_data_log_force[2204] <= 16'h0000;
      coeffs_in_data_log_force[2205] <= 16'h0000;
      coeffs_in_data_log_force[2206] <= 16'h0000;
      coeffs_in_data_log_force[2207] <= 16'h0000;
      coeffs_in_data_log_force[2208] <= 16'h0000;
      coeffs_in_data_log_force[2209] <= 16'h0000;
      coeffs_in_data_log_force[2210] <= 16'h0000;
      coeffs_in_data_log_force[2211] <= 16'h0000;
      coeffs_in_data_log_force[2212] <= 16'h0000;
      coeffs_in_data_log_force[2213] <= 16'h0000;
      coeffs_in_data_log_force[2214] <= 16'h0000;
      coeffs_in_data_log_force[2215] <= 16'h0000;
      coeffs_in_data_log_force[2216] <= 16'h0000;
      coeffs_in_data_log_force[2217] <= 16'h0000;
      coeffs_in_data_log_force[2218] <= 16'h0000;
      coeffs_in_data_log_force[2219] <= 16'h0000;
      coeffs_in_data_log_force[2220] <= 16'h0000;
      coeffs_in_data_log_force[2221] <= 16'h0000;
      coeffs_in_data_log_force[2222] <= 16'h0000;
      coeffs_in_data_log_force[2223] <= 16'h0000;
      coeffs_in_data_log_force[2224] <= 16'h0000;
      coeffs_in_data_log_force[2225] <= 16'h0000;
      coeffs_in_data_log_force[2226] <= 16'h0000;
      coeffs_in_data_log_force[2227] <= 16'h0000;
      coeffs_in_data_log_force[2228] <= 16'h0000;
      coeffs_in_data_log_force[2229] <= 16'h0000;
      coeffs_in_data_log_force[2230] <= 16'h0000;
      coeffs_in_data_log_force[2231] <= 16'h0000;
      coeffs_in_data_log_force[2232] <= 16'h0000;
      coeffs_in_data_log_force[2233] <= 16'h0000;
      coeffs_in_data_log_force[2234] <= 16'h0000;
      coeffs_in_data_log_force[2235] <= 16'h0000;
      coeffs_in_data_log_force[2236] <= 16'h0000;
      coeffs_in_data_log_force[2237] <= 16'h0000;
      coeffs_in_data_log_force[2238] <= 16'h0000;
      coeffs_in_data_log_force[2239] <= 16'h0000;
      coeffs_in_data_log_force[2240] <= 16'h0000;
      coeffs_in_data_log_force[2241] <= 16'h0000;
      coeffs_in_data_log_force[2242] <= 16'h0000;
      coeffs_in_data_log_force[2243] <= 16'h0000;
      coeffs_in_data_log_force[2244] <= 16'h0000;
      coeffs_in_data_log_force[2245] <= 16'h0000;
      coeffs_in_data_log_force[2246] <= 16'h0000;
      coeffs_in_data_log_force[2247] <= 16'h0000;
      coeffs_in_data_log_force[2248] <= 16'h0000;
      coeffs_in_data_log_force[2249] <= 16'h0000;
      coeffs_in_data_log_force[2250] <= 16'h0000;
      coeffs_in_data_log_force[2251] <= 16'h0000;
      coeffs_in_data_log_force[2252] <= 16'h0000;
      coeffs_in_data_log_force[2253] <= 16'h0000;
      coeffs_in_data_log_force[2254] <= 16'h0000;
      coeffs_in_data_log_force[2255] <= 16'h0000;
      coeffs_in_data_log_force[2256] <= 16'h0000;
      coeffs_in_data_log_force[2257] <= 16'h0000;
      coeffs_in_data_log_force[2258] <= 16'h0000;
      coeffs_in_data_log_force[2259] <= 16'h0000;
      coeffs_in_data_log_force[2260] <= 16'h0000;
      coeffs_in_data_log_force[2261] <= 16'h0000;
      coeffs_in_data_log_force[2262] <= 16'h0000;
      coeffs_in_data_log_force[2263] <= 16'h0000;
      coeffs_in_data_log_force[2264] <= 16'h0000;
      coeffs_in_data_log_force[2265] <= 16'h0000;
      coeffs_in_data_log_force[2266] <= 16'h0000;
      coeffs_in_data_log_force[2267] <= 16'h0000;
      coeffs_in_data_log_force[2268] <= 16'h0000;
      coeffs_in_data_log_force[2269] <= 16'h0000;
      coeffs_in_data_log_force[2270] <= 16'h0000;
      coeffs_in_data_log_force[2271] <= 16'h0000;
      coeffs_in_data_log_force[2272] <= 16'h0000;
      coeffs_in_data_log_force[2273] <= 16'h0000;
      coeffs_in_data_log_force[2274] <= 16'h0000;
      coeffs_in_data_log_force[2275] <= 16'h0000;
      coeffs_in_data_log_force[2276] <= 16'h0000;
      coeffs_in_data_log_force[2277] <= 16'h0000;
      coeffs_in_data_log_force[2278] <= 16'h0000;
      coeffs_in_data_log_force[2279] <= 16'h0000;
      coeffs_in_data_log_force[2280] <= 16'h0000;
      coeffs_in_data_log_force[2281] <= 16'h0000;
      coeffs_in_data_log_force[2282] <= 16'h0000;
      coeffs_in_data_log_force[2283] <= 16'h0000;
      coeffs_in_data_log_force[2284] <= 16'h0000;
      coeffs_in_data_log_force[2285] <= 16'h0000;
      coeffs_in_data_log_force[2286] <= 16'h0000;
      coeffs_in_data_log_force[2287] <= 16'h0000;
      coeffs_in_data_log_force[2288] <= 16'h0000;
      coeffs_in_data_log_force[2289] <= 16'h0000;
      coeffs_in_data_log_force[2290] <= 16'h0000;
      coeffs_in_data_log_force[2291] <= 16'h0000;
      coeffs_in_data_log_force[2292] <= 16'h0000;
      coeffs_in_data_log_force[2293] <= 16'h0000;
      coeffs_in_data_log_force[2294] <= 16'h0000;
      coeffs_in_data_log_force[2295] <= 16'h0000;
      coeffs_in_data_log_force[2296] <= 16'h0000;
      coeffs_in_data_log_force[2297] <= 16'h0000;
      coeffs_in_data_log_force[2298] <= 16'h0000;
      coeffs_in_data_log_force[2299] <= 16'h0000;
      coeffs_in_data_log_force[2300] <= 16'h0000;
      coeffs_in_data_log_force[2301] <= 16'h0000;
      coeffs_in_data_log_force[2302] <= 16'h0000;
      coeffs_in_data_log_force[2303] <= 16'h0000;
      coeffs_in_data_log_force[2304] <= 16'h0000;
      coeffs_in_data_log_force[2305] <= 16'h0000;
      coeffs_in_data_log_force[2306] <= 16'h0000;
      coeffs_in_data_log_force[2307] <= 16'h0000;
      coeffs_in_data_log_force[2308] <= 16'h0000;
      coeffs_in_data_log_force[2309] <= 16'h0000;
      coeffs_in_data_log_force[2310] <= 16'h0000;
      coeffs_in_data_log_force[2311] <= 16'h0000;
      coeffs_in_data_log_force[2312] <= 16'h0000;
      coeffs_in_data_log_force[2313] <= 16'h0000;
      coeffs_in_data_log_force[2314] <= 16'h0000;
      coeffs_in_data_log_force[2315] <= 16'h0000;
      coeffs_in_data_log_force[2316] <= 16'h0000;
      coeffs_in_data_log_force[2317] <= 16'h0000;
      coeffs_in_data_log_force[2318] <= 16'h0000;
      coeffs_in_data_log_force[2319] <= 16'h0000;
      coeffs_in_data_log_force[2320] <= 16'h0000;
      coeffs_in_data_log_force[2321] <= 16'h0000;
      coeffs_in_data_log_force[2322] <= 16'h0000;
      coeffs_in_data_log_force[2323] <= 16'h0000;
      coeffs_in_data_log_force[2324] <= 16'h0000;
      coeffs_in_data_log_force[2325] <= 16'h0000;
      coeffs_in_data_log_force[2326] <= 16'h0000;
      coeffs_in_data_log_force[2327] <= 16'h0000;
      coeffs_in_data_log_force[2328] <= 16'h0000;
      coeffs_in_data_log_force[2329] <= 16'h0000;
      coeffs_in_data_log_force[2330] <= 16'h0000;
      coeffs_in_data_log_force[2331] <= 16'h0000;
      coeffs_in_data_log_force[2332] <= 16'h0000;
      coeffs_in_data_log_force[2333] <= 16'h0000;
      coeffs_in_data_log_force[2334] <= 16'h0000;
      coeffs_in_data_log_force[2335] <= 16'h0000;
      coeffs_in_data_log_force[2336] <= 16'h0000;
      coeffs_in_data_log_force[2337] <= 16'h0000;
      coeffs_in_data_log_force[2338] <= 16'h0000;
      coeffs_in_data_log_force[2339] <= 16'h0000;
      coeffs_in_data_log_force[2340] <= 16'h0000;
      coeffs_in_data_log_force[2341] <= 16'h0000;
      coeffs_in_data_log_force[2342] <= 16'h0000;
      coeffs_in_data_log_force[2343] <= 16'h0000;
      coeffs_in_data_log_force[2344] <= 16'h0000;
      coeffs_in_data_log_force[2345] <= 16'h0000;
      coeffs_in_data_log_force[2346] <= 16'h0000;
      coeffs_in_data_log_force[2347] <= 16'h0000;
      coeffs_in_data_log_force[2348] <= 16'h0000;
      coeffs_in_data_log_force[2349] <= 16'h0000;
      coeffs_in_data_log_force[2350] <= 16'h0000;
      coeffs_in_data_log_force[2351] <= 16'h0000;
      coeffs_in_data_log_force[2352] <= 16'h0000;
      coeffs_in_data_log_force[2353] <= 16'h0000;
      coeffs_in_data_log_force[2354] <= 16'h0000;
      coeffs_in_data_log_force[2355] <= 16'h0000;
      coeffs_in_data_log_force[2356] <= 16'h0000;
      coeffs_in_data_log_force[2357] <= 16'h0000;
      coeffs_in_data_log_force[2358] <= 16'h0000;
      coeffs_in_data_log_force[2359] <= 16'h0000;
      coeffs_in_data_log_force[2360] <= 16'h0000;
      coeffs_in_data_log_force[2361] <= 16'h0000;
      coeffs_in_data_log_force[2362] <= 16'h0000;
      coeffs_in_data_log_force[2363] <= 16'h0000;
      coeffs_in_data_log_force[2364] <= 16'h0000;
      coeffs_in_data_log_force[2365] <= 16'h0000;
      coeffs_in_data_log_force[2366] <= 16'h0000;
      coeffs_in_data_log_force[2367] <= 16'h0000;
      coeffs_in_data_log_force[2368] <= 16'h0000;
      coeffs_in_data_log_force[2369] <= 16'h0000;
      coeffs_in_data_log_force[2370] <= 16'h0000;
      coeffs_in_data_log_force[2371] <= 16'h0000;
      coeffs_in_data_log_force[2372] <= 16'h0000;
      coeffs_in_data_log_force[2373] <= 16'h0000;
      coeffs_in_data_log_force[2374] <= 16'h0000;
      coeffs_in_data_log_force[2375] <= 16'h0000;
      coeffs_in_data_log_force[2376] <= 16'h0000;
      coeffs_in_data_log_force[2377] <= 16'h0000;
      coeffs_in_data_log_force[2378] <= 16'h0000;
      coeffs_in_data_log_force[2379] <= 16'h0000;
      coeffs_in_data_log_force[2380] <= 16'h0000;
      coeffs_in_data_log_force[2381] <= 16'h0000;
      coeffs_in_data_log_force[2382] <= 16'h0000;
      coeffs_in_data_log_force[2383] <= 16'h0000;
      coeffs_in_data_log_force[2384] <= 16'h0000;
      coeffs_in_data_log_force[2385] <= 16'h0000;
      coeffs_in_data_log_force[2386] <= 16'h0000;
      coeffs_in_data_log_force[2387] <= 16'h0000;
      coeffs_in_data_log_force[2388] <= 16'h0000;
      coeffs_in_data_log_force[2389] <= 16'h0000;
      coeffs_in_data_log_force[2390] <= 16'h0000;
      coeffs_in_data_log_force[2391] <= 16'h0000;
      coeffs_in_data_log_force[2392] <= 16'h0000;
      coeffs_in_data_log_force[2393] <= 16'h0000;
      coeffs_in_data_log_force[2394] <= 16'h0000;
      coeffs_in_data_log_force[2395] <= 16'h0000;
      coeffs_in_data_log_force[2396] <= 16'h0000;
      coeffs_in_data_log_force[2397] <= 16'h0000;
      coeffs_in_data_log_force[2398] <= 16'h0000;
      coeffs_in_data_log_force[2399] <= 16'h0000;
      coeffs_in_data_log_force[2400] <= 16'h0000;
      coeffs_in_data_log_force[2401] <= 16'h0000;
      coeffs_in_data_log_force[2402] <= 16'h0000;
      coeffs_in_data_log_force[2403] <= 16'h0000;
      coeffs_in_data_log_force[2404] <= 16'h0000;
      coeffs_in_data_log_force[2405] <= 16'h0000;
      coeffs_in_data_log_force[2406] <= 16'h0000;
      coeffs_in_data_log_force[2407] <= 16'h0000;
      coeffs_in_data_log_force[2408] <= 16'h0000;
      coeffs_in_data_log_force[2409] <= 16'h0000;
      coeffs_in_data_log_force[2410] <= 16'h0000;
      coeffs_in_data_log_force[2411] <= 16'h0000;
      coeffs_in_data_log_force[2412] <= 16'h0000;
      coeffs_in_data_log_force[2413] <= 16'h0000;
      coeffs_in_data_log_force[2414] <= 16'h0000;
      coeffs_in_data_log_force[2415] <= 16'h0000;
      coeffs_in_data_log_force[2416] <= 16'h0000;
      coeffs_in_data_log_force[2417] <= 16'h0000;
      coeffs_in_data_log_force[2418] <= 16'h0000;
      coeffs_in_data_log_force[2419] <= 16'h0000;
      coeffs_in_data_log_force[2420] <= 16'h0000;
      coeffs_in_data_log_force[2421] <= 16'h0000;
      coeffs_in_data_log_force[2422] <= 16'h0000;
      coeffs_in_data_log_force[2423] <= 16'h0000;
      coeffs_in_data_log_force[2424] <= 16'h0000;
      coeffs_in_data_log_force[2425] <= 16'h0000;
      coeffs_in_data_log_force[2426] <= 16'h0000;
      coeffs_in_data_log_force[2427] <= 16'h0000;
      coeffs_in_data_log_force[2428] <= 16'h0000;
      coeffs_in_data_log_force[2429] <= 16'h0000;
      coeffs_in_data_log_force[2430] <= 16'h0000;
      coeffs_in_data_log_force[2431] <= 16'h0000;
      coeffs_in_data_log_force[2432] <= 16'h0000;
      coeffs_in_data_log_force[2433] <= 16'h0000;
      coeffs_in_data_log_force[2434] <= 16'h0000;
      coeffs_in_data_log_force[2435] <= 16'h0000;
      coeffs_in_data_log_force[2436] <= 16'h0000;
      coeffs_in_data_log_force[2437] <= 16'h0000;
      coeffs_in_data_log_force[2438] <= 16'h0000;
      coeffs_in_data_log_force[2439] <= 16'h0000;
      coeffs_in_data_log_force[2440] <= 16'h0000;
      coeffs_in_data_log_force[2441] <= 16'h0000;
      coeffs_in_data_log_force[2442] <= 16'h0000;
      coeffs_in_data_log_force[2443] <= 16'h0000;
      coeffs_in_data_log_force[2444] <= 16'h0000;
      coeffs_in_data_log_force[2445] <= 16'h0000;
      coeffs_in_data_log_force[2446] <= 16'h0000;
      coeffs_in_data_log_force[2447] <= 16'h0000;
      coeffs_in_data_log_force[2448] <= 16'h0000;
      coeffs_in_data_log_force[2449] <= 16'h0000;
      coeffs_in_data_log_force[2450] <= 16'h0000;
      coeffs_in_data_log_force[2451] <= 16'h0000;
      coeffs_in_data_log_force[2452] <= 16'h0000;
      coeffs_in_data_log_force[2453] <= 16'h0000;
      coeffs_in_data_log_force[2454] <= 16'h0000;
      coeffs_in_data_log_force[2455] <= 16'h0000;
      coeffs_in_data_log_force[2456] <= 16'h0000;
      coeffs_in_data_log_force[2457] <= 16'h0000;
      coeffs_in_data_log_force[2458] <= 16'h0000;
      coeffs_in_data_log_force[2459] <= 16'h0000;
      coeffs_in_data_log_force[2460] <= 16'h0000;
      coeffs_in_data_log_force[2461] <= 16'h0000;
      coeffs_in_data_log_force[2462] <= 16'h0000;
      coeffs_in_data_log_force[2463] <= 16'h0000;
      coeffs_in_data_log_force[2464] <= 16'h0000;
      coeffs_in_data_log_force[2465] <= 16'h0000;
      coeffs_in_data_log_force[2466] <= 16'h0000;
      coeffs_in_data_log_force[2467] <= 16'h0000;
      coeffs_in_data_log_force[2468] <= 16'h0000;
      coeffs_in_data_log_force[2469] <= 16'h0000;
      coeffs_in_data_log_force[2470] <= 16'h0000;
      coeffs_in_data_log_force[2471] <= 16'h0000;
      coeffs_in_data_log_force[2472] <= 16'h0000;
      coeffs_in_data_log_force[2473] <= 16'h0000;
      coeffs_in_data_log_force[2474] <= 16'h0000;
      coeffs_in_data_log_force[2475] <= 16'h0000;
      coeffs_in_data_log_force[2476] <= 16'h0000;
      coeffs_in_data_log_force[2477] <= 16'h0000;
      coeffs_in_data_log_force[2478] <= 16'h0000;
      coeffs_in_data_log_force[2479] <= 16'h0000;
      coeffs_in_data_log_force[2480] <= 16'h0000;
      coeffs_in_data_log_force[2481] <= 16'h0000;
      coeffs_in_data_log_force[2482] <= 16'h0000;
      coeffs_in_data_log_force[2483] <= 16'h0000;
      coeffs_in_data_log_force[2484] <= 16'h0000;
      coeffs_in_data_log_force[2485] <= 16'h0000;
      coeffs_in_data_log_force[2486] <= 16'h0000;
      coeffs_in_data_log_force[2487] <= 16'h0000;
      coeffs_in_data_log_force[2488] <= 16'h0000;
      coeffs_in_data_log_force[2489] <= 16'h0000;
      coeffs_in_data_log_force[2490] <= 16'h0000;
      coeffs_in_data_log_force[2491] <= 16'h0000;
      coeffs_in_data_log_force[2492] <= 16'h0000;
      coeffs_in_data_log_force[2493] <= 16'h0000;
      coeffs_in_data_log_force[2494] <= 16'h0000;
      coeffs_in_data_log_force[2495] <= 16'h0000;
      coeffs_in_data_log_force[2496] <= 16'h0000;
      coeffs_in_data_log_force[2497] <= 16'h0000;
      coeffs_in_data_log_force[2498] <= 16'h0000;
      coeffs_in_data_log_force[2499] <= 16'h0000;
      coeffs_in_data_log_force[2500] <= 16'h0000;
      coeffs_in_data_log_force[2501] <= 16'h0000;
      coeffs_in_data_log_force[2502] <= 16'h0000;
      coeffs_in_data_log_force[2503] <= 16'h0000;
      coeffs_in_data_log_force[2504] <= 16'h0000;
      coeffs_in_data_log_force[2505] <= 16'h0000;
      coeffs_in_data_log_force[2506] <= 16'h0000;
      coeffs_in_data_log_force[2507] <= 16'h0000;
      coeffs_in_data_log_force[2508] <= 16'h0000;
      coeffs_in_data_log_force[2509] <= 16'h0000;
      coeffs_in_data_log_force[2510] <= 16'h0000;
      coeffs_in_data_log_force[2511] <= 16'h0000;
      coeffs_in_data_log_force[2512] <= 16'h0000;
      coeffs_in_data_log_force[2513] <= 16'h0000;
      coeffs_in_data_log_force[2514] <= 16'h0000;
      coeffs_in_data_log_force[2515] <= 16'h0000;
      coeffs_in_data_log_force[2516] <= 16'h0000;
      coeffs_in_data_log_force[2517] <= 16'h0000;
      coeffs_in_data_log_force[2518] <= 16'h0000;
      coeffs_in_data_log_force[2519] <= 16'h0000;
      coeffs_in_data_log_force[2520] <= 16'h0000;
      coeffs_in_data_log_force[2521] <= 16'h0000;
      coeffs_in_data_log_force[2522] <= 16'h0000;
      coeffs_in_data_log_force[2523] <= 16'h0000;
      coeffs_in_data_log_force[2524] <= 16'h0000;
      coeffs_in_data_log_force[2525] <= 16'h0000;
      coeffs_in_data_log_force[2526] <= 16'h0000;
      coeffs_in_data_log_force[2527] <= 16'h0000;
      coeffs_in_data_log_force[2528] <= 16'h0000;
      coeffs_in_data_log_force[2529] <= 16'h0000;
      coeffs_in_data_log_force[2530] <= 16'h0000;
      coeffs_in_data_log_force[2531] <= 16'h0000;
      coeffs_in_data_log_force[2532] <= 16'h0000;
      coeffs_in_data_log_force[2533] <= 16'h0000;
      coeffs_in_data_log_force[2534] <= 16'h0000;
      coeffs_in_data_log_force[2535] <= 16'h0000;
      coeffs_in_data_log_force[2536] <= 16'h0000;
      coeffs_in_data_log_force[2537] <= 16'h0000;
      coeffs_in_data_log_force[2538] <= 16'h0000;
      coeffs_in_data_log_force[2539] <= 16'h0000;
      coeffs_in_data_log_force[2540] <= 16'h0000;
      coeffs_in_data_log_force[2541] <= 16'h0000;
      coeffs_in_data_log_force[2542] <= 16'h0000;
      coeffs_in_data_log_force[2543] <= 16'h0000;
      coeffs_in_data_log_force[2544] <= 16'h0000;
      coeffs_in_data_log_force[2545] <= 16'h0000;
      coeffs_in_data_log_force[2546] <= 16'h0000;
      coeffs_in_data_log_force[2547] <= 16'h0000;
      coeffs_in_data_log_force[2548] <= 16'h0000;
      coeffs_in_data_log_force[2549] <= 16'h0000;
      coeffs_in_data_log_force[2550] <= 16'h0000;
      coeffs_in_data_log_force[2551] <= 16'h0000;
      coeffs_in_data_log_force[2552] <= 16'h0000;
      coeffs_in_data_log_force[2553] <= 16'h0000;
      coeffs_in_data_log_force[2554] <= 16'h0000;
      coeffs_in_data_log_force[2555] <= 16'h0000;
      coeffs_in_data_log_force[2556] <= 16'h0000;
      coeffs_in_data_log_force[2557] <= 16'h0000;
      coeffs_in_data_log_force[2558] <= 16'h0000;
      coeffs_in_data_log_force[2559] <= 16'h0000;
      coeffs_in_data_log_force[2560] <= 16'h0000;
      coeffs_in_data_log_force[2561] <= 16'h0000;
      coeffs_in_data_log_force[2562] <= 16'h0000;
      coeffs_in_data_log_force[2563] <= 16'h0000;
      coeffs_in_data_log_force[2564] <= 16'h0000;
      coeffs_in_data_log_force[2565] <= 16'h0000;
      coeffs_in_data_log_force[2566] <= 16'h0000;
      coeffs_in_data_log_force[2567] <= 16'h0000;
      coeffs_in_data_log_force[2568] <= 16'h0000;
      coeffs_in_data_log_force[2569] <= 16'h0000;
      coeffs_in_data_log_force[2570] <= 16'h0000;
      coeffs_in_data_log_force[2571] <= 16'h0000;
      coeffs_in_data_log_force[2572] <= 16'h0000;
      coeffs_in_data_log_force[2573] <= 16'h0000;
      coeffs_in_data_log_force[2574] <= 16'h0000;
      coeffs_in_data_log_force[2575] <= 16'h0000;
      coeffs_in_data_log_force[2576] <= 16'h0000;
      coeffs_in_data_log_force[2577] <= 16'h0000;
      coeffs_in_data_log_force[2578] <= 16'h0000;
      coeffs_in_data_log_force[2579] <= 16'h0000;
      coeffs_in_data_log_force[2580] <= 16'h0000;
      coeffs_in_data_log_force[2581] <= 16'h0000;
      coeffs_in_data_log_force[2582] <= 16'h0000;
      coeffs_in_data_log_force[2583] <= 16'h0000;
      coeffs_in_data_log_force[2584] <= 16'h0000;
      coeffs_in_data_log_force[2585] <= 16'h0000;
      coeffs_in_data_log_force[2586] <= 16'h0000;
      coeffs_in_data_log_force[2587] <= 16'h0000;
      coeffs_in_data_log_force[2588] <= 16'h0000;
      coeffs_in_data_log_force[2589] <= 16'h0000;
      coeffs_in_data_log_force[2590] <= 16'h0000;
      coeffs_in_data_log_force[2591] <= 16'h0000;
      coeffs_in_data_log_force[2592] <= 16'h0000;
      coeffs_in_data_log_force[2593] <= 16'h0000;
      coeffs_in_data_log_force[2594] <= 16'h0000;
      coeffs_in_data_log_force[2595] <= 16'h0000;
      coeffs_in_data_log_force[2596] <= 16'h0000;
      coeffs_in_data_log_force[2597] <= 16'h0000;
      coeffs_in_data_log_force[2598] <= 16'h0000;
      coeffs_in_data_log_force[2599] <= 16'h0000;
      coeffs_in_data_log_force[2600] <= 16'h0000;
      coeffs_in_data_log_force[2601] <= 16'h0000;
      coeffs_in_data_log_force[2602] <= 16'h0000;
      coeffs_in_data_log_force[2603] <= 16'h0000;
      coeffs_in_data_log_force[2604] <= 16'h0000;
      coeffs_in_data_log_force[2605] <= 16'h0000;
      coeffs_in_data_log_force[2606] <= 16'h0000;
      coeffs_in_data_log_force[2607] <= 16'h0000;
      coeffs_in_data_log_force[2608] <= 16'h0000;
      coeffs_in_data_log_force[2609] <= 16'h0000;
      coeffs_in_data_log_force[2610] <= 16'h0000;
      coeffs_in_data_log_force[2611] <= 16'h0000;
      coeffs_in_data_log_force[2612] <= 16'h0000;
      coeffs_in_data_log_force[2613] <= 16'h0000;
      coeffs_in_data_log_force[2614] <= 16'h0000;
      coeffs_in_data_log_force[2615] <= 16'h0000;
      coeffs_in_data_log_force[2616] <= 16'h0000;
      coeffs_in_data_log_force[2617] <= 16'h0000;
      coeffs_in_data_log_force[2618] <= 16'h0000;
      coeffs_in_data_log_force[2619] <= 16'h0000;
      coeffs_in_data_log_force[2620] <= 16'h0000;
      coeffs_in_data_log_force[2621] <= 16'h0000;
      coeffs_in_data_log_force[2622] <= 16'h0000;
      coeffs_in_data_log_force[2623] <= 16'h0000;
      coeffs_in_data_log_force[2624] <= 16'h0000;
      coeffs_in_data_log_force[2625] <= 16'h0000;
      coeffs_in_data_log_force[2626] <= 16'h0000;
      coeffs_in_data_log_force[2627] <= 16'h0000;
      coeffs_in_data_log_force[2628] <= 16'h0000;
      coeffs_in_data_log_force[2629] <= 16'h0000;
      coeffs_in_data_log_force[2630] <= 16'h0000;
      coeffs_in_data_log_force[2631] <= 16'h0000;
      coeffs_in_data_log_force[2632] <= 16'h0000;
      coeffs_in_data_log_force[2633] <= 16'h0000;
      coeffs_in_data_log_force[2634] <= 16'h0000;
      coeffs_in_data_log_force[2635] <= 16'h0000;
      coeffs_in_data_log_force[2636] <= 16'h0000;
      coeffs_in_data_log_force[2637] <= 16'h0000;
      coeffs_in_data_log_force[2638] <= 16'h0000;
      coeffs_in_data_log_force[2639] <= 16'h0000;
      coeffs_in_data_log_force[2640] <= 16'h0000;
      coeffs_in_data_log_force[2641] <= 16'h0000;
      coeffs_in_data_log_force[2642] <= 16'h0000;
      coeffs_in_data_log_force[2643] <= 16'h0000;
      coeffs_in_data_log_force[2644] <= 16'h0000;
      coeffs_in_data_log_force[2645] <= 16'h0000;
      coeffs_in_data_log_force[2646] <= 16'h0000;
      coeffs_in_data_log_force[2647] <= 16'h0000;
      coeffs_in_data_log_force[2648] <= 16'h0000;
      coeffs_in_data_log_force[2649] <= 16'h0000;
      coeffs_in_data_log_force[2650] <= 16'h0000;
      coeffs_in_data_log_force[2651] <= 16'h0000;
      coeffs_in_data_log_force[2652] <= 16'h0000;
      coeffs_in_data_log_force[2653] <= 16'h0000;
      coeffs_in_data_log_force[2654] <= 16'h0000;
      coeffs_in_data_log_force[2655] <= 16'h0000;
      coeffs_in_data_log_force[2656] <= 16'h0000;
      coeffs_in_data_log_force[2657] <= 16'h0000;
      coeffs_in_data_log_force[2658] <= 16'h0000;
      coeffs_in_data_log_force[2659] <= 16'h0000;
      coeffs_in_data_log_force[2660] <= 16'h0000;
      coeffs_in_data_log_force[2661] <= 16'h0000;
      coeffs_in_data_log_force[2662] <= 16'h0000;
      coeffs_in_data_log_force[2663] <= 16'h0000;
      coeffs_in_data_log_force[2664] <= 16'h0000;
      coeffs_in_data_log_force[2665] <= 16'h0000;
      coeffs_in_data_log_force[2666] <= 16'h0000;
      coeffs_in_data_log_force[2667] <= 16'h0000;
      coeffs_in_data_log_force[2668] <= 16'h0000;
      coeffs_in_data_log_force[2669] <= 16'h0000;
      coeffs_in_data_log_force[2670] <= 16'h0000;
      coeffs_in_data_log_force[2671] <= 16'h0000;
      coeffs_in_data_log_force[2672] <= 16'h0000;
      coeffs_in_data_log_force[2673] <= 16'h0000;
      coeffs_in_data_log_force[2674] <= 16'h0000;
      coeffs_in_data_log_force[2675] <= 16'h0000;
      coeffs_in_data_log_force[2676] <= 16'h0000;
      coeffs_in_data_log_force[2677] <= 16'h0000;
      coeffs_in_data_log_force[2678] <= 16'h0000;
      coeffs_in_data_log_force[2679] <= 16'h0000;
      coeffs_in_data_log_force[2680] <= 16'h0000;
      coeffs_in_data_log_force[2681] <= 16'h0000;
      coeffs_in_data_log_force[2682] <= 16'h0000;
      coeffs_in_data_log_force[2683] <= 16'h0000;
      coeffs_in_data_log_force[2684] <= 16'h0000;
      coeffs_in_data_log_force[2685] <= 16'h0000;
      coeffs_in_data_log_force[2686] <= 16'h0000;
      coeffs_in_data_log_force[2687] <= 16'h0000;
      coeffs_in_data_log_force[2688] <= 16'h0000;
      coeffs_in_data_log_force[2689] <= 16'h0000;
      coeffs_in_data_log_force[2690] <= 16'h0000;
      coeffs_in_data_log_force[2691] <= 16'h0000;
      coeffs_in_data_log_force[2692] <= 16'h0000;
      coeffs_in_data_log_force[2693] <= 16'h0000;
      coeffs_in_data_log_force[2694] <= 16'h0000;
      coeffs_in_data_log_force[2695] <= 16'h0000;
      coeffs_in_data_log_force[2696] <= 16'h0000;
      coeffs_in_data_log_force[2697] <= 16'h0000;
      coeffs_in_data_log_force[2698] <= 16'h0000;
      coeffs_in_data_log_force[2699] <= 16'h0000;
      coeffs_in_data_log_force[2700] <= 16'h0000;
      coeffs_in_data_log_force[2701] <= 16'h0000;
      coeffs_in_data_log_force[2702] <= 16'h0000;
      coeffs_in_data_log_force[2703] <= 16'h0000;
      coeffs_in_data_log_force[2704] <= 16'h0000;
      coeffs_in_data_log_force[2705] <= 16'h0000;
      coeffs_in_data_log_force[2706] <= 16'h0000;
      coeffs_in_data_log_force[2707] <= 16'h0000;
      coeffs_in_data_log_force[2708] <= 16'h0000;
      coeffs_in_data_log_force[2709] <= 16'h0000;
      coeffs_in_data_log_force[2710] <= 16'h0000;
      coeffs_in_data_log_force[2711] <= 16'h0000;
      coeffs_in_data_log_force[2712] <= 16'h0000;
      coeffs_in_data_log_force[2713] <= 16'h0000;
      coeffs_in_data_log_force[2714] <= 16'h0000;
      coeffs_in_data_log_force[2715] <= 16'h0000;
      coeffs_in_data_log_force[2716] <= 16'h0000;
      coeffs_in_data_log_force[2717] <= 16'h0000;
      coeffs_in_data_log_force[2718] <= 16'h0000;
      coeffs_in_data_log_force[2719] <= 16'h0000;
      coeffs_in_data_log_force[2720] <= 16'h0000;
      coeffs_in_data_log_force[2721] <= 16'h0000;
      coeffs_in_data_log_force[2722] <= 16'h0000;
      coeffs_in_data_log_force[2723] <= 16'h0000;
      coeffs_in_data_log_force[2724] <= 16'h0000;
      coeffs_in_data_log_force[2725] <= 16'h0000;
      coeffs_in_data_log_force[2726] <= 16'h0000;
      coeffs_in_data_log_force[2727] <= 16'h0000;
      coeffs_in_data_log_force[2728] <= 16'h0000;
      coeffs_in_data_log_force[2729] <= 16'h0000;
      coeffs_in_data_log_force[2730] <= 16'h0000;
      coeffs_in_data_log_force[2731] <= 16'h0000;
      coeffs_in_data_log_force[2732] <= 16'h0000;
      coeffs_in_data_log_force[2733] <= 16'h0000;
      coeffs_in_data_log_force[2734] <= 16'h0000;
      coeffs_in_data_log_force[2735] <= 16'h0000;
      coeffs_in_data_log_force[2736] <= 16'h0000;
      coeffs_in_data_log_force[2737] <= 16'h0000;
      coeffs_in_data_log_force[2738] <= 16'h0000;
      coeffs_in_data_log_force[2739] <= 16'h0000;
      coeffs_in_data_log_force[2740] <= 16'h0000;
      coeffs_in_data_log_force[2741] <= 16'h0000;
      coeffs_in_data_log_force[2742] <= 16'h0000;
      coeffs_in_data_log_force[2743] <= 16'h0000;
      coeffs_in_data_log_force[2744] <= 16'h0000;
      coeffs_in_data_log_force[2745] <= 16'h0000;
      coeffs_in_data_log_force[2746] <= 16'h0000;
      coeffs_in_data_log_force[2747] <= 16'h0000;
      coeffs_in_data_log_force[2748] <= 16'h0000;
      coeffs_in_data_log_force[2749] <= 16'h0000;
      coeffs_in_data_log_force[2750] <= 16'h0000;
      coeffs_in_data_log_force[2751] <= 16'h0000;
      coeffs_in_data_log_force[2752] <= 16'h0000;
      coeffs_in_data_log_force[2753] <= 16'h0000;
      coeffs_in_data_log_force[2754] <= 16'h0000;
      coeffs_in_data_log_force[2755] <= 16'h0000;
      coeffs_in_data_log_force[2756] <= 16'h0000;
      coeffs_in_data_log_force[2757] <= 16'h0000;
      coeffs_in_data_log_force[2758] <= 16'h0000;
      coeffs_in_data_log_force[2759] <= 16'h0000;
      coeffs_in_data_log_force[2760] <= 16'h0000;
      coeffs_in_data_log_force[2761] <= 16'h0000;
      coeffs_in_data_log_force[2762] <= 16'h0000;
      coeffs_in_data_log_force[2763] <= 16'h0000;
      coeffs_in_data_log_force[2764] <= 16'h0000;
      coeffs_in_data_log_force[2765] <= 16'h0000;
      coeffs_in_data_log_force[2766] <= 16'h0000;
      coeffs_in_data_log_force[2767] <= 16'h0000;
      coeffs_in_data_log_force[2768] <= 16'h0000;
      coeffs_in_data_log_force[2769] <= 16'h0000;
      coeffs_in_data_log_force[2770] <= 16'h0000;
      coeffs_in_data_log_force[2771] <= 16'h0000;
      coeffs_in_data_log_force[2772] <= 16'h0000;
      coeffs_in_data_log_force[2773] <= 16'h0000;
      coeffs_in_data_log_force[2774] <= 16'h0000;
      coeffs_in_data_log_force[2775] <= 16'h0000;
      coeffs_in_data_log_force[2776] <= 16'h0000;
      coeffs_in_data_log_force[2777] <= 16'h0000;
      coeffs_in_data_log_force[2778] <= 16'h0000;
      coeffs_in_data_log_force[2779] <= 16'h0000;
      coeffs_in_data_log_force[2780] <= 16'h0000;
      coeffs_in_data_log_force[2781] <= 16'h0000;
      coeffs_in_data_log_force[2782] <= 16'h0000;
      coeffs_in_data_log_force[2783] <= 16'h0000;
      coeffs_in_data_log_force[2784] <= 16'h0000;
      coeffs_in_data_log_force[2785] <= 16'h0000;
      coeffs_in_data_log_force[2786] <= 16'h0000;
      coeffs_in_data_log_force[2787] <= 16'h0000;
      coeffs_in_data_log_force[2788] <= 16'h0000;
      coeffs_in_data_log_force[2789] <= 16'h0000;
      coeffs_in_data_log_force[2790] <= 16'h0000;
      coeffs_in_data_log_force[2791] <= 16'h0000;
      coeffs_in_data_log_force[2792] <= 16'h0000;
      coeffs_in_data_log_force[2793] <= 16'h0000;
      coeffs_in_data_log_force[2794] <= 16'h0000;
      coeffs_in_data_log_force[2795] <= 16'h0000;
      coeffs_in_data_log_force[2796] <= 16'h0000;
      coeffs_in_data_log_force[2797] <= 16'h0000;
      coeffs_in_data_log_force[2798] <= 16'h0000;
      coeffs_in_data_log_force[2799] <= 16'h0000;
      coeffs_in_data_log_force[2800] <= 16'h0000;
      coeffs_in_data_log_force[2801] <= 16'h0000;
      coeffs_in_data_log_force[2802] <= 16'h0000;
      coeffs_in_data_log_force[2803] <= 16'h0000;
      coeffs_in_data_log_force[2804] <= 16'h0000;
      coeffs_in_data_log_force[2805] <= 16'h0000;
      coeffs_in_data_log_force[2806] <= 16'h0000;
      coeffs_in_data_log_force[2807] <= 16'h0000;
      coeffs_in_data_log_force[2808] <= 16'h0000;
      coeffs_in_data_log_force[2809] <= 16'h0000;
      coeffs_in_data_log_force[2810] <= 16'h0000;
      coeffs_in_data_log_force[2811] <= 16'h0000;
      coeffs_in_data_log_force[2812] <= 16'h0000;
      coeffs_in_data_log_force[2813] <= 16'h0000;
      coeffs_in_data_log_force[2814] <= 16'h0000;
      coeffs_in_data_log_force[2815] <= 16'h0000;
      coeffs_in_data_log_force[2816] <= 16'h0000;
      coeffs_in_data_log_force[2817] <= 16'h0000;
      coeffs_in_data_log_force[2818] <= 16'h0000;
      coeffs_in_data_log_force[2819] <= 16'h0000;
      coeffs_in_data_log_force[2820] <= 16'h0000;
      coeffs_in_data_log_force[2821] <= 16'h0000;
      coeffs_in_data_log_force[2822] <= 16'h0000;
      coeffs_in_data_log_force[2823] <= 16'h0000;
      coeffs_in_data_log_force[2824] <= 16'h0000;
      coeffs_in_data_log_force[2825] <= 16'h0000;
      coeffs_in_data_log_force[2826] <= 16'h0000;
      coeffs_in_data_log_force[2827] <= 16'h0000;
      coeffs_in_data_log_force[2828] <= 16'h0000;
      coeffs_in_data_log_force[2829] <= 16'h0000;
      coeffs_in_data_log_force[2830] <= 16'h0000;
      coeffs_in_data_log_force[2831] <= 16'h0000;
      coeffs_in_data_log_force[2832] <= 16'h0000;
      coeffs_in_data_log_force[2833] <= 16'h0000;
      coeffs_in_data_log_force[2834] <= 16'h0000;
      coeffs_in_data_log_force[2835] <= 16'h0000;
      coeffs_in_data_log_force[2836] <= 16'h0000;
      coeffs_in_data_log_force[2837] <= 16'h0000;
      coeffs_in_data_log_force[2838] <= 16'h0000;
      coeffs_in_data_log_force[2839] <= 16'h0000;
      coeffs_in_data_log_force[2840] <= 16'h0000;
      coeffs_in_data_log_force[2841] <= 16'h0000;
      coeffs_in_data_log_force[2842] <= 16'h0000;
      coeffs_in_data_log_force[2843] <= 16'h0000;
      coeffs_in_data_log_force[2844] <= 16'h0000;
      coeffs_in_data_log_force[2845] <= 16'h0000;
      coeffs_in_data_log_force[2846] <= 16'h0000;
      coeffs_in_data_log_force[2847] <= 16'h0000;
      coeffs_in_data_log_force[2848] <= 16'h0000;
      coeffs_in_data_log_force[2849] <= 16'h0000;
      coeffs_in_data_log_force[2850] <= 16'h0000;
      coeffs_in_data_log_force[2851] <= 16'h0000;
      coeffs_in_data_log_force[2852] <= 16'h0000;
      coeffs_in_data_log_force[2853] <= 16'h0000;
      coeffs_in_data_log_force[2854] <= 16'h0000;
      coeffs_in_data_log_force[2855] <= 16'h0000;
      coeffs_in_data_log_force[2856] <= 16'h0000;
      coeffs_in_data_log_force[2857] <= 16'h0000;
      coeffs_in_data_log_force[2858] <= 16'h0000;
      coeffs_in_data_log_force[2859] <= 16'h0000;
      coeffs_in_data_log_force[2860] <= 16'h0000;
      coeffs_in_data_log_force[2861] <= 16'h0000;
      coeffs_in_data_log_force[2862] <= 16'h0000;
      coeffs_in_data_log_force[2863] <= 16'h0000;
      coeffs_in_data_log_force[2864] <= 16'h0000;
      coeffs_in_data_log_force[2865] <= 16'h0000;
      coeffs_in_data_log_force[2866] <= 16'h0000;
      coeffs_in_data_log_force[2867] <= 16'h0000;
      coeffs_in_data_log_force[2868] <= 16'h0000;
      coeffs_in_data_log_force[2869] <= 16'h0000;
      coeffs_in_data_log_force[2870] <= 16'h0000;
      coeffs_in_data_log_force[2871] <= 16'h0000;
      coeffs_in_data_log_force[2872] <= 16'h0000;
      coeffs_in_data_log_force[2873] <= 16'h0000;
      coeffs_in_data_log_force[2874] <= 16'h0000;
      coeffs_in_data_log_force[2875] <= 16'h0000;
      coeffs_in_data_log_force[2876] <= 16'h0000;
      coeffs_in_data_log_force[2877] <= 16'h0000;
      coeffs_in_data_log_force[2878] <= 16'h0000;
      coeffs_in_data_log_force[2879] <= 16'h0000;
      coeffs_in_data_log_force[2880] <= 16'h0000;
      coeffs_in_data_log_force[2881] <= 16'h0000;
      coeffs_in_data_log_force[2882] <= 16'h0000;
      coeffs_in_data_log_force[2883] <= 16'h0000;
      coeffs_in_data_log_force[2884] <= 16'h0000;
      coeffs_in_data_log_force[2885] <= 16'h0000;
      coeffs_in_data_log_force[2886] <= 16'h0000;
      coeffs_in_data_log_force[2887] <= 16'h0000;
      coeffs_in_data_log_force[2888] <= 16'h0000;
      coeffs_in_data_log_force[2889] <= 16'h0000;
      coeffs_in_data_log_force[2890] <= 16'h0000;
      coeffs_in_data_log_force[2891] <= 16'h0000;
      coeffs_in_data_log_force[2892] <= 16'h0000;
      coeffs_in_data_log_force[2893] <= 16'h0000;
      coeffs_in_data_log_force[2894] <= 16'h0000;
      coeffs_in_data_log_force[2895] <= 16'h0000;
      coeffs_in_data_log_force[2896] <= 16'h0000;
      coeffs_in_data_log_force[2897] <= 16'h0000;
      coeffs_in_data_log_force[2898] <= 16'h0000;
      coeffs_in_data_log_force[2899] <= 16'h0000;
      coeffs_in_data_log_force[2900] <= 16'h0000;
      coeffs_in_data_log_force[2901] <= 16'h0000;
      coeffs_in_data_log_force[2902] <= 16'h0000;
      coeffs_in_data_log_force[2903] <= 16'h0000;
      coeffs_in_data_log_force[2904] <= 16'h0000;
      coeffs_in_data_log_force[2905] <= 16'h0000;
      coeffs_in_data_log_force[2906] <= 16'h0000;
      coeffs_in_data_log_force[2907] <= 16'h0000;
      coeffs_in_data_log_force[2908] <= 16'h0000;
      coeffs_in_data_log_force[2909] <= 16'h0000;
      coeffs_in_data_log_force[2910] <= 16'h0000;
      coeffs_in_data_log_force[2911] <= 16'h0000;
      coeffs_in_data_log_force[2912] <= 16'h0000;
      coeffs_in_data_log_force[2913] <= 16'h0000;
      coeffs_in_data_log_force[2914] <= 16'h0000;
      coeffs_in_data_log_force[2915] <= 16'h0000;
      coeffs_in_data_log_force[2916] <= 16'h0000;
      coeffs_in_data_log_force[2917] <= 16'h0000;
      coeffs_in_data_log_force[2918] <= 16'h0000;
      coeffs_in_data_log_force[2919] <= 16'h0000;
      coeffs_in_data_log_force[2920] <= 16'h0000;
      coeffs_in_data_log_force[2921] <= 16'h0000;
      coeffs_in_data_log_force[2922] <= 16'h0000;
      coeffs_in_data_log_force[2923] <= 16'h0000;
      coeffs_in_data_log_force[2924] <= 16'h0000;
      coeffs_in_data_log_force[2925] <= 16'h0000;
      coeffs_in_data_log_force[2926] <= 16'h0000;
      coeffs_in_data_log_force[2927] <= 16'h0000;
      coeffs_in_data_log_force[2928] <= 16'h0000;
      coeffs_in_data_log_force[2929] <= 16'h0000;
      coeffs_in_data_log_force[2930] <= 16'h0000;
      coeffs_in_data_log_force[2931] <= 16'h0000;
      coeffs_in_data_log_force[2932] <= 16'h0000;
      coeffs_in_data_log_force[2933] <= 16'h0000;
      coeffs_in_data_log_force[2934] <= 16'h0000;
      coeffs_in_data_log_force[2935] <= 16'h0000;
      coeffs_in_data_log_force[2936] <= 16'h0000;
      coeffs_in_data_log_force[2937] <= 16'h0000;
      coeffs_in_data_log_force[2938] <= 16'h0000;
      coeffs_in_data_log_force[2939] <= 16'h0000;
      coeffs_in_data_log_force[2940] <= 16'h0000;
      coeffs_in_data_log_force[2941] <= 16'h0000;
      coeffs_in_data_log_force[2942] <= 16'h0000;
      coeffs_in_data_log_force[2943] <= 16'h0000;
      coeffs_in_data_log_force[2944] <= 16'h0000;
      coeffs_in_data_log_force[2945] <= 16'h0000;
      coeffs_in_data_log_force[2946] <= 16'h0000;
      coeffs_in_data_log_force[2947] <= 16'h0000;
      coeffs_in_data_log_force[2948] <= 16'h0000;
      coeffs_in_data_log_force[2949] <= 16'h0000;
      coeffs_in_data_log_force[2950] <= 16'h0000;
      coeffs_in_data_log_force[2951] <= 16'h0000;
      coeffs_in_data_log_force[2952] <= 16'h0000;
      coeffs_in_data_log_force[2953] <= 16'h0000;
      coeffs_in_data_log_force[2954] <= 16'h0000;
      coeffs_in_data_log_force[2955] <= 16'h0000;
      coeffs_in_data_log_force[2956] <= 16'h0000;
      coeffs_in_data_log_force[2957] <= 16'h0000;
      coeffs_in_data_log_force[2958] <= 16'h0000;
      coeffs_in_data_log_force[2959] <= 16'h0000;
      coeffs_in_data_log_force[2960] <= 16'h0000;
      coeffs_in_data_log_force[2961] <= 16'h0000;
      coeffs_in_data_log_force[2962] <= 16'h0000;
      coeffs_in_data_log_force[2963] <= 16'h0000;
      coeffs_in_data_log_force[2964] <= 16'h0000;
      coeffs_in_data_log_force[2965] <= 16'h0000;
      coeffs_in_data_log_force[2966] <= 16'h0000;
      coeffs_in_data_log_force[2967] <= 16'h0000;
      coeffs_in_data_log_force[2968] <= 16'h0000;
      coeffs_in_data_log_force[2969] <= 16'h0000;
      coeffs_in_data_log_force[2970] <= 16'h0000;
      coeffs_in_data_log_force[2971] <= 16'h0000;
      coeffs_in_data_log_force[2972] <= 16'h0000;
      coeffs_in_data_log_force[2973] <= 16'h0000;
      coeffs_in_data_log_force[2974] <= 16'h0000;
      coeffs_in_data_log_force[2975] <= 16'h0000;
      coeffs_in_data_log_force[2976] <= 16'h0000;
      coeffs_in_data_log_force[2977] <= 16'h0000;
      coeffs_in_data_log_force[2978] <= 16'h0000;
      coeffs_in_data_log_force[2979] <= 16'h0000;
      coeffs_in_data_log_force[2980] <= 16'h0000;
      coeffs_in_data_log_force[2981] <= 16'h0000;
      coeffs_in_data_log_force[2982] <= 16'h0000;
      coeffs_in_data_log_force[2983] <= 16'h0000;
      coeffs_in_data_log_force[2984] <= 16'h0000;
      coeffs_in_data_log_force[2985] <= 16'h0000;
      coeffs_in_data_log_force[2986] <= 16'h0000;
      coeffs_in_data_log_force[2987] <= 16'h0000;
      coeffs_in_data_log_force[2988] <= 16'h0000;
      coeffs_in_data_log_force[2989] <= 16'h0000;
      coeffs_in_data_log_force[2990] <= 16'h0000;
      coeffs_in_data_log_force[2991] <= 16'h0000;
      coeffs_in_data_log_force[2992] <= 16'h0000;
      coeffs_in_data_log_force[2993] <= 16'h0000;
      coeffs_in_data_log_force[2994] <= 16'h0000;
      coeffs_in_data_log_force[2995] <= 16'h0000;
      coeffs_in_data_log_force[2996] <= 16'h0000;
      coeffs_in_data_log_force[2997] <= 16'h0000;
      coeffs_in_data_log_force[2998] <= 16'h0000;
      coeffs_in_data_log_force[2999] <= 16'h0000;
      coeffs_in_data_log_force[3000] <= 16'h0000;
      coeffs_in_data_log_force[3001] <= 16'h0000;
      coeffs_in_data_log_force[3002] <= 16'h0000;
      coeffs_in_data_log_force[3003] <= 16'h0000;
      coeffs_in_data_log_force[3004] <= 16'h0000;
      coeffs_in_data_log_force[3005] <= 16'h0000;
      coeffs_in_data_log_force[3006] <= 16'h0000;
      coeffs_in_data_log_force[3007] <= 16'h0000;
      coeffs_in_data_log_force[3008] <= 16'h0000;
      coeffs_in_data_log_force[3009] <= 16'h0000;
      coeffs_in_data_log_force[3010] <= 16'h0000;
      coeffs_in_data_log_force[3011] <= 16'h0000;
      coeffs_in_data_log_force[3012] <= 16'h0000;
      coeffs_in_data_log_force[3013] <= 16'h0000;
      coeffs_in_data_log_force[3014] <= 16'h0000;
      coeffs_in_data_log_force[3015] <= 16'h0000;
      coeffs_in_data_log_force[3016] <= 16'h0000;
      coeffs_in_data_log_force[3017] <= 16'h0000;
      coeffs_in_data_log_force[3018] <= 16'h0000;
      coeffs_in_data_log_force[3019] <= 16'h0000;
      coeffs_in_data_log_force[3020] <= 16'h0000;
      coeffs_in_data_log_force[3021] <= 16'h0000;
      coeffs_in_data_log_force[3022] <= 16'h0000;
      coeffs_in_data_log_force[3023] <= 16'h0000;
      coeffs_in_data_log_force[3024] <= 16'h0000;
      coeffs_in_data_log_force[3025] <= 16'h0000;
      coeffs_in_data_log_force[3026] <= 16'h0000;
      coeffs_in_data_log_force[3027] <= 16'h0000;
      coeffs_in_data_log_force[3028] <= 16'h0000;
      coeffs_in_data_log_force[3029] <= 16'h0000;
      coeffs_in_data_log_force[3030] <= 16'h0000;
      coeffs_in_data_log_force[3031] <= 16'h0000;
      coeffs_in_data_log_force[3032] <= 16'h0000;
      coeffs_in_data_log_force[3033] <= 16'h0000;
      coeffs_in_data_log_force[3034] <= 16'h0000;
      coeffs_in_data_log_force[3035] <= 16'h0000;
      coeffs_in_data_log_force[3036] <= 16'h0000;
      coeffs_in_data_log_force[3037] <= 16'h0000;
      coeffs_in_data_log_force[3038] <= 16'h0000;
      coeffs_in_data_log_force[3039] <= 16'h0000;
      coeffs_in_data_log_force[3040] <= 16'h0000;
      coeffs_in_data_log_force[3041] <= 16'h0000;
      coeffs_in_data_log_force[3042] <= 16'h0000;
      coeffs_in_data_log_force[3043] <= 16'h0000;
      coeffs_in_data_log_force[3044] <= 16'h0000;
      coeffs_in_data_log_force[3045] <= 16'h0000;
      coeffs_in_data_log_force[3046] <= 16'h0000;
      coeffs_in_data_log_force[3047] <= 16'h0000;
      coeffs_in_data_log_force[3048] <= 16'h0000;
      coeffs_in_data_log_force[3049] <= 16'h0000;
      coeffs_in_data_log_force[3050] <= 16'h0000;
      coeffs_in_data_log_force[3051] <= 16'h0000;
      coeffs_in_data_log_force[3052] <= 16'h0000;
      coeffs_in_data_log_force[3053] <= 16'h0000;
      coeffs_in_data_log_force[3054] <= 16'h0000;
      coeffs_in_data_log_force[3055] <= 16'h0000;
      coeffs_in_data_log_force[3056] <= 16'h0000;
      coeffs_in_data_log_force[3057] <= 16'h0000;
      coeffs_in_data_log_force[3058] <= 16'h0000;
      coeffs_in_data_log_force[3059] <= 16'h0000;
      coeffs_in_data_log_force[3060] <= 16'h0000;
      coeffs_in_data_log_force[3061] <= 16'h0000;
      coeffs_in_data_log_force[3062] <= 16'h0000;
      coeffs_in_data_log_force[3063] <= 16'h0000;
      coeffs_in_data_log_force[3064] <= 16'h0000;
      coeffs_in_data_log_force[3065] <= 16'h0000;
      coeffs_in_data_log_force[3066] <= 16'h0000;
      coeffs_in_data_log_force[3067] <= 16'h0000;
      coeffs_in_data_log_force[3068] <= 16'h0000;
      coeffs_in_data_log_force[3069] <= 16'h0000;
      coeffs_in_data_log_force[3070] <= 16'h0000;
      coeffs_in_data_log_force[3071] <= 16'h0000;
      coeffs_in_data_log_force[3072] <= 16'h0000;
      coeffs_in_data_log_force[3073] <= 16'h0000;
      coeffs_in_data_log_force[3074] <= 16'h0000;
      coeffs_in_data_log_force[3075] <= 16'h0000;
      coeffs_in_data_log_force[3076] <= 16'h0000;
      coeffs_in_data_log_force[3077] <= 16'h0000;
      coeffs_in_data_log_force[3078] <= 16'h0000;
      coeffs_in_data_log_force[3079] <= 16'h0000;
      coeffs_in_data_log_force[3080] <= 16'h0000;
      coeffs_in_data_log_force[3081] <= 16'h0000;
      coeffs_in_data_log_force[3082] <= 16'h0000;
      coeffs_in_data_log_force[3083] <= 16'h0000;
      coeffs_in_data_log_force[3084] <= 16'h0000;
      coeffs_in_data_log_force[3085] <= 16'h0000;
      coeffs_in_data_log_force[3086] <= 16'h0000;
      coeffs_in_data_log_force[3087] <= 16'h0000;
      coeffs_in_data_log_force[3088] <= 16'h0000;
      coeffs_in_data_log_force[3089] <= 16'h0000;
      coeffs_in_data_log_force[3090] <= 16'h0000;
      coeffs_in_data_log_force[3091] <= 16'h0000;
      coeffs_in_data_log_force[3092] <= 16'h0000;
      coeffs_in_data_log_force[3093] <= 16'h0000;
      coeffs_in_data_log_force[3094] <= 16'h0000;
      coeffs_in_data_log_force[3095] <= 16'h0000;
      coeffs_in_data_log_force[3096] <= 16'h0000;
      coeffs_in_data_log_force[3097] <= 16'h0000;
      coeffs_in_data_log_force[3098] <= 16'h0000;
      coeffs_in_data_log_force[3099] <= 16'h0000;
      coeffs_in_data_log_force[3100] <= 16'h0000;
      coeffs_in_data_log_force[3101] <= 16'h0000;
      coeffs_in_data_log_force[3102] <= 16'h0000;
      coeffs_in_data_log_force[3103] <= 16'h0000;
      coeffs_in_data_log_force[3104] <= 16'h0000;
      coeffs_in_data_log_force[3105] <= 16'h0000;
      coeffs_in_data_log_force[3106] <= 16'h0000;
      coeffs_in_data_log_force[3107] <= 16'h0000;
      coeffs_in_data_log_force[3108] <= 16'h0000;
      coeffs_in_data_log_force[3109] <= 16'h0000;
      coeffs_in_data_log_force[3110] <= 16'h0000;
      coeffs_in_data_log_force[3111] <= 16'h0000;
      coeffs_in_data_log_force[3112] <= 16'h0000;
      coeffs_in_data_log_force[3113] <= 16'h0000;
      coeffs_in_data_log_force[3114] <= 16'h0000;
      coeffs_in_data_log_force[3115] <= 16'h0000;
      coeffs_in_data_log_force[3116] <= 16'h0000;
      coeffs_in_data_log_force[3117] <= 16'h0000;
      coeffs_in_data_log_force[3118] <= 16'h0000;
      coeffs_in_data_log_force[3119] <= 16'h0000;
      coeffs_in_data_log_force[3120] <= 16'h0000;
      coeffs_in_data_log_force[3121] <= 16'h0000;
      coeffs_in_data_log_force[3122] <= 16'h0000;
      coeffs_in_data_log_force[3123] <= 16'h0000;
      coeffs_in_data_log_force[3124] <= 16'h0000;
      coeffs_in_data_log_force[3125] <= 16'h0000;
      coeffs_in_data_log_force[3126] <= 16'h0000;
      coeffs_in_data_log_force[3127] <= 16'h0000;
      coeffs_in_data_log_force[3128] <= 16'h0000;
      coeffs_in_data_log_force[3129] <= 16'h0000;
      coeffs_in_data_log_force[3130] <= 16'h0000;
      coeffs_in_data_log_force[3131] <= 16'h0000;
      coeffs_in_data_log_force[3132] <= 16'h0000;
      coeffs_in_data_log_force[3133] <= 16'h0000;
      coeffs_in_data_log_force[3134] <= 16'h0000;
      coeffs_in_data_log_force[3135] <= 16'h0000;
      coeffs_in_data_log_force[3136] <= 16'h0000;
      coeffs_in_data_log_force[3137] <= 16'h0000;
      coeffs_in_data_log_force[3138] <= 16'h0000;
      coeffs_in_data_log_force[3139] <= 16'h0000;
      coeffs_in_data_log_force[3140] <= 16'h0000;
      coeffs_in_data_log_force[3141] <= 16'h0000;
      coeffs_in_data_log_force[3142] <= 16'h0000;
      coeffs_in_data_log_force[3143] <= 16'h0000;
      coeffs_in_data_log_force[3144] <= 16'h0000;
      coeffs_in_data_log_force[3145] <= 16'h0000;
      coeffs_in_data_log_force[3146] <= 16'h0000;
      coeffs_in_data_log_force[3147] <= 16'h0000;
      coeffs_in_data_log_force[3148] <= 16'h0000;
      coeffs_in_data_log_force[3149] <= 16'h0000;
      coeffs_in_data_log_force[3150] <= 16'h0000;
      coeffs_in_data_log_force[3151] <= 16'h0000;
      coeffs_in_data_log_force[3152] <= 16'h0000;
      coeffs_in_data_log_force[3153] <= 16'h0000;
      coeffs_in_data_log_force[3154] <= 16'h0000;
      coeffs_in_data_log_force[3155] <= 16'h0000;
      coeffs_in_data_log_force[3156] <= 16'h0000;
      coeffs_in_data_log_force[3157] <= 16'h0000;
      coeffs_in_data_log_force[3158] <= 16'h0000;
      coeffs_in_data_log_force[3159] <= 16'h0000;
      coeffs_in_data_log_force[3160] <= 16'h0000;
      coeffs_in_data_log_force[3161] <= 16'h0000;
      coeffs_in_data_log_force[3162] <= 16'h0000;
      coeffs_in_data_log_force[3163] <= 16'h0000;
      coeffs_in_data_log_force[3164] <= 16'h0000;
      coeffs_in_data_log_force[3165] <= 16'h0000;
      coeffs_in_data_log_force[3166] <= 16'h0000;
      coeffs_in_data_log_force[3167] <= 16'h0000;
      coeffs_in_data_log_force[3168] <= 16'h0000;
      coeffs_in_data_log_force[3169] <= 16'h0000;
      coeffs_in_data_log_force[3170] <= 16'h0000;
      coeffs_in_data_log_force[3171] <= 16'h0000;
      coeffs_in_data_log_force[3172] <= 16'h0000;
      coeffs_in_data_log_force[3173] <= 16'h0000;
      coeffs_in_data_log_force[3174] <= 16'h0000;
      coeffs_in_data_log_force[3175] <= 16'h0000;
      coeffs_in_data_log_force[3176] <= 16'h0000;
      coeffs_in_data_log_force[3177] <= 16'h0000;
      coeffs_in_data_log_force[3178] <= 16'h0000;
      coeffs_in_data_log_force[3179] <= 16'h0000;
      coeffs_in_data_log_force[3180] <= 16'h0000;
      coeffs_in_data_log_force[3181] <= 16'h0000;
      coeffs_in_data_log_force[3182] <= 16'h0000;
      coeffs_in_data_log_force[3183] <= 16'h0000;
      coeffs_in_data_log_force[3184] <= 16'h0000;
      coeffs_in_data_log_force[3185] <= 16'h0000;
      coeffs_in_data_log_force[3186] <= 16'h0000;
      coeffs_in_data_log_force[3187] <= 16'h0000;
      coeffs_in_data_log_force[3188] <= 16'h0000;
      coeffs_in_data_log_force[3189] <= 16'h0000;
      coeffs_in_data_log_force[3190] <= 16'h0000;
      coeffs_in_data_log_force[3191] <= 16'h0000;
      coeffs_in_data_log_force[3192] <= 16'h0000;
      coeffs_in_data_log_force[3193] <= 16'h0000;
      coeffs_in_data_log_force[3194] <= 16'h0000;
      coeffs_in_data_log_force[3195] <= 16'h0000;
      coeffs_in_data_log_force[3196] <= 16'h0000;
      coeffs_in_data_log_force[3197] <= 16'h0000;
      coeffs_in_data_log_force[3198] <= 16'h0000;
      coeffs_in_data_log_force[3199] <= 16'h0000;
      coeffs_in_data_log_force[3200] <= 16'h0000;
      coeffs_in_data_log_force[3201] <= 16'h0000;
      coeffs_in_data_log_force[3202] <= 16'h0000;
      coeffs_in_data_log_force[3203] <= 16'h0000;
      coeffs_in_data_log_force[3204] <= 16'h0000;
      coeffs_in_data_log_force[3205] <= 16'h0000;
      coeffs_in_data_log_force[3206] <= 16'h0000;
      coeffs_in_data_log_force[3207] <= 16'h0000;
      coeffs_in_data_log_force[3208] <= 16'h0000;
      coeffs_in_data_log_force[3209] <= 16'h0000;
      coeffs_in_data_log_force[3210] <= 16'h0000;
      coeffs_in_data_log_force[3211] <= 16'h0000;
      coeffs_in_data_log_force[3212] <= 16'h0000;
      coeffs_in_data_log_force[3213] <= 16'h0000;
      coeffs_in_data_log_force[3214] <= 16'h0000;
      coeffs_in_data_log_force[3215] <= 16'h0000;
      coeffs_in_data_log_force[3216] <= 16'h0000;
      coeffs_in_data_log_force[3217] <= 16'h0000;
      coeffs_in_data_log_force[3218] <= 16'h0000;
      coeffs_in_data_log_force[3219] <= 16'h0000;
      coeffs_in_data_log_force[3220] <= 16'h0000;
      coeffs_in_data_log_force[3221] <= 16'h0000;
      coeffs_in_data_log_force[3222] <= 16'h0000;
      coeffs_in_data_log_force[3223] <= 16'h0000;
      coeffs_in_data_log_force[3224] <= 16'h0000;
      coeffs_in_data_log_force[3225] <= 16'h0000;
      coeffs_in_data_log_force[3226] <= 16'h0000;
      coeffs_in_data_log_force[3227] <= 16'h0000;
      coeffs_in_data_log_force[3228] <= 16'h0000;
      coeffs_in_data_log_force[3229] <= 16'h0000;
      coeffs_in_data_log_force[3230] <= 16'h0000;
      coeffs_in_data_log_force[3231] <= 16'h0000;
      coeffs_in_data_log_force[3232] <= 16'h0000;
      coeffs_in_data_log_force[3233] <= 16'h0000;
      coeffs_in_data_log_force[3234] <= 16'h0000;
      coeffs_in_data_log_force[3235] <= 16'h0000;
      coeffs_in_data_log_force[3236] <= 16'h0000;
      coeffs_in_data_log_force[3237] <= 16'h0000;
      coeffs_in_data_log_force[3238] <= 16'h0000;
      coeffs_in_data_log_force[3239] <= 16'h0000;
      coeffs_in_data_log_force[3240] <= 16'h0000;
      coeffs_in_data_log_force[3241] <= 16'h0000;
      coeffs_in_data_log_force[3242] <= 16'h0000;
      coeffs_in_data_log_force[3243] <= 16'h0000;
      coeffs_in_data_log_force[3244] <= 16'h0000;
      coeffs_in_data_log_force[3245] <= 16'h0000;
      coeffs_in_data_log_force[3246] <= 16'h0000;
      coeffs_in_data_log_force[3247] <= 16'h0000;
      coeffs_in_data_log_force[3248] <= 16'h0000;
      coeffs_in_data_log_force[3249] <= 16'h0000;
      coeffs_in_data_log_force[3250] <= 16'h0000;
      coeffs_in_data_log_force[3251] <= 16'h0000;
      coeffs_in_data_log_force[3252] <= 16'h0000;
      coeffs_in_data_log_force[3253] <= 16'h0000;
      coeffs_in_data_log_force[3254] <= 16'h0000;
      coeffs_in_data_log_force[3255] <= 16'h0000;
      coeffs_in_data_log_force[3256] <= 16'h0000;
      coeffs_in_data_log_force[3257] <= 16'h0000;
      coeffs_in_data_log_force[3258] <= 16'h0000;
      coeffs_in_data_log_force[3259] <= 16'h0000;
      coeffs_in_data_log_force[3260] <= 16'h0000;
      coeffs_in_data_log_force[3261] <= 16'h0000;
      coeffs_in_data_log_force[3262] <= 16'h0000;
      coeffs_in_data_log_force[3263] <= 16'h0000;
      coeffs_in_data_log_force[3264] <= 16'h0000;
      coeffs_in_data_log_force[3265] <= 16'h0000;
      coeffs_in_data_log_force[3266] <= 16'h0000;
      coeffs_in_data_log_force[3267] <= 16'h0000;
      coeffs_in_data_log_force[3268] <= 16'h0000;
      coeffs_in_data_log_force[3269] <= 16'h0000;
      coeffs_in_data_log_force[3270] <= 16'h0000;
      coeffs_in_data_log_force[3271] <= 16'h0000;
      coeffs_in_data_log_force[3272] <= 16'h0000;
      coeffs_in_data_log_force[3273] <= 16'h0000;
      coeffs_in_data_log_force[3274] <= 16'h0000;
      coeffs_in_data_log_force[3275] <= 16'h0000;
      coeffs_in_data_log_force[3276] <= 16'h0000;
      coeffs_in_data_log_force[3277] <= 16'h0000;
      coeffs_in_data_log_force[3278] <= 16'h0000;
      coeffs_in_data_log_force[3279] <= 16'h0000;
      coeffs_in_data_log_force[3280] <= 16'h0000;
      coeffs_in_data_log_force[3281] <= 16'h0000;
      coeffs_in_data_log_force[3282] <= 16'h0000;
      coeffs_in_data_log_force[3283] <= 16'h0000;
      coeffs_in_data_log_force[3284] <= 16'h0000;
      coeffs_in_data_log_force[3285] <= 16'h0000;
      coeffs_in_data_log_force[3286] <= 16'h0000;
      coeffs_in_data_log_force[3287] <= 16'h0000;
      coeffs_in_data_log_force[3288] <= 16'h0000;
      coeffs_in_data_log_force[3289] <= 16'h0000;
      coeffs_in_data_log_force[3290] <= 16'h0000;
      coeffs_in_data_log_force[3291] <= 16'h0000;
      coeffs_in_data_log_force[3292] <= 16'h0000;
      coeffs_in_data_log_force[3293] <= 16'h0000;
      coeffs_in_data_log_force[3294] <= 16'h0000;
      coeffs_in_data_log_force[3295] <= 16'h0000;
      coeffs_in_data_log_force[3296] <= 16'h0000;
      coeffs_in_data_log_force[3297] <= 16'h0000;
      coeffs_in_data_log_force[3298] <= 16'h0000;
      coeffs_in_data_log_force[3299] <= 16'h0000;
      coeffs_in_data_log_force[3300] <= 16'h0000;
      coeffs_in_data_log_force[3301] <= 16'h0000;
      coeffs_in_data_log_force[3302] <= 16'h0000;
      coeffs_in_data_log_force[3303] <= 16'h0000;
      coeffs_in_data_log_force[3304] <= 16'h0000;
      coeffs_in_data_log_force[3305] <= 16'h0000;
      coeffs_in_data_log_force[3306] <= 16'h0000;
      coeffs_in_data_log_force[3307] <= 16'h0000;
      coeffs_in_data_log_force[3308] <= 16'h0000;
      coeffs_in_data_log_force[3309] <= 16'h0000;
      coeffs_in_data_log_force[3310] <= 16'h0000;
      coeffs_in_data_log_force[3311] <= 16'h0000;
      coeffs_in_data_log_force[3312] <= 16'h0000;
      coeffs_in_data_log_force[3313] <= 16'h0000;
      coeffs_in_data_log_force[3314] <= 16'h0000;
      coeffs_in_data_log_force[3315] <= 16'h0000;
      coeffs_in_data_log_force[3316] <= 16'h0000;
      coeffs_in_data_log_force[3317] <= 16'h0000;
      coeffs_in_data_log_force[3318] <= 16'h0000;
      coeffs_in_data_log_force[3319] <= 16'h0000;
      coeffs_in_data_log_force[3320] <= 16'h0000;
      coeffs_in_data_log_force[3321] <= 16'h0000;
      coeffs_in_data_log_force[3322] <= 16'h0000;
      coeffs_in_data_log_force[3323] <= 16'h0000;
      coeffs_in_data_log_force[3324] <= 16'h0000;
      coeffs_in_data_log_force[3325] <= 16'h0000;
      coeffs_in_data_log_force[3326] <= 16'h0000;
      coeffs_in_data_log_force[3327] <= 16'h0000;
      coeffs_in_data_log_force[3328] <= 16'h0000;
      coeffs_in_data_log_force[3329] <= 16'h0000;
      coeffs_in_data_log_force[3330] <= 16'h0000;
      coeffs_in_data_log_force[3331] <= 16'h0000;
      coeffs_in_data_log_force[3332] <= 16'h0000;
      coeffs_in_data_log_force[3333] <= 16'h0000;
      coeffs_in_data_log_force[3334] <= 16'h0000;
      coeffs_in_data_log_force[3335] <= 16'h0000;
      coeffs_in_data_log_force[3336] <= 16'h0000;
      coeffs_in_data_log_force[3337] <= 16'h0000;
      coeffs_in_data_log_force[3338] <= 16'h0000;
      coeffs_in_data_log_force[3339] <= 16'h0000;
      coeffs_in_data_log_force[3340] <= 16'h0000;
      coeffs_in_data_log_force[3341] <= 16'h0000;
      coeffs_in_data_log_force[3342] <= 16'h0000;
      coeffs_in_data_log_force[3343] <= 16'h0000;
      coeffs_in_data_log_force[3344] <= 16'h0000;
      coeffs_in_data_log_force[3345] <= 16'h0000;
      coeffs_in_data_log_force[3346] <= 16'h0000;
      coeffs_in_data_log_force[3347] <= 16'h0000;
      coeffs_in_data_log_force[3348] <= 16'h0000;
      coeffs_in_data_log_force[3349] <= 16'h0000;
      coeffs_in_data_log_force[3350] <= 16'h0000;
      coeffs_in_data_log_force[3351] <= 16'h0000;
      coeffs_in_data_log_force[3352] <= 16'h0000;
      coeffs_in_data_log_force[3353] <= 16'h0000;
      coeffs_in_data_log_force[3354] <= 16'h0000;
      coeffs_in_data_log_force[3355] <= 16'h0000;
      coeffs_in_data_log_force[3356] <= 16'h0000;
      coeffs_in_data_log_force[3357] <= 16'h0000;
      coeffs_in_data_log_force[3358] <= 16'h0000;
      coeffs_in_data_log_force[3359] <= 16'h0000;
      coeffs_in_data_log_force[3360] <= 16'h0000;
      coeffs_in_data_log_force[3361] <= 16'h0000;
      coeffs_in_data_log_force[3362] <= 16'h0000;
      coeffs_in_data_log_force[3363] <= 16'h0000;
      coeffs_in_data_log_force[3364] <= 16'h0000;
      coeffs_in_data_log_force[3365] <= 16'h0000;
      coeffs_in_data_log_force[3366] <= 16'h0000;
      coeffs_in_data_log_force[3367] <= 16'h0000;
      coeffs_in_data_log_force[3368] <= 16'h0000;
      coeffs_in_data_log_force[3369] <= 16'h0000;
      coeffs_in_data_log_force[3370] <= 16'h0000;
      coeffs_in_data_log_force[3371] <= 16'h0000;
      coeffs_in_data_log_force[3372] <= 16'h0000;
      coeffs_in_data_log_force[3373] <= 16'h0000;
      coeffs_in_data_log_force[3374] <= 16'h0000;
      coeffs_in_data_log_force[3375] <= 16'h0000;
      coeffs_in_data_log_force[3376] <= 16'h0000;
      coeffs_in_data_log_force[3377] <= 16'h0000;
      coeffs_in_data_log_force[3378] <= 16'h0000;
      coeffs_in_data_log_force[3379] <= 16'h0000;
      coeffs_in_data_log_force[3380] <= 16'h0000;
      coeffs_in_data_log_force[3381] <= 16'h0000;
      coeffs_in_data_log_force[3382] <= 16'h0000;
      coeffs_in_data_log_force[3383] <= 16'h0000;
      coeffs_in_data_log_force[3384] <= 16'h0000;
      coeffs_in_data_log_force[3385] <= 16'h0000;
      coeffs_in_data_log_force[3386] <= 16'h0000;
      coeffs_in_data_log_force[3387] <= 16'h0000;
      coeffs_in_data_log_force[3388] <= 16'h0000;
      coeffs_in_data_log_force[3389] <= 16'h0000;
      coeffs_in_data_log_force[3390] <= 16'h0000;
      coeffs_in_data_log_force[3391] <= 16'h0000;
      coeffs_in_data_log_force[3392] <= 16'h0000;
      coeffs_in_data_log_force[3393] <= 16'h0000;
      coeffs_in_data_log_force[3394] <= 16'h0000;
      coeffs_in_data_log_force[3395] <= 16'h0000;
      coeffs_in_data_log_force[3396] <= 16'h0000;
      coeffs_in_data_log_force[3397] <= 16'h0000;
      coeffs_in_data_log_force[3398] <= 16'h0000;
      coeffs_in_data_log_force[3399] <= 16'h0000;
      coeffs_in_data_log_force[3400] <= 16'h0000;
      coeffs_in_data_log_force[3401] <= 16'h0000;
      coeffs_in_data_log_force[3402] <= 16'h0000;
      coeffs_in_data_log_force[3403] <= 16'h0000;
      coeffs_in_data_log_force[3404] <= 16'h0000;
      coeffs_in_data_log_force[3405] <= 16'h0000;
      coeffs_in_data_log_force[3406] <= 16'h0000;
      coeffs_in_data_log_force[3407] <= 16'h0000;
      coeffs_in_data_log_force[3408] <= 16'h0000;
      coeffs_in_data_log_force[3409] <= 16'h0000;
      coeffs_in_data_log_force[3410] <= 16'h0000;
      coeffs_in_data_log_force[3411] <= 16'h0000;
      coeffs_in_data_log_force[3412] <= 16'h0000;
      coeffs_in_data_log_force[3413] <= 16'h0000;
      coeffs_in_data_log_force[3414] <= 16'h0000;
      coeffs_in_data_log_force[3415] <= 16'h0000;
      coeffs_in_data_log_force[3416] <= 16'h0000;
      coeffs_in_data_log_force[3417] <= 16'h0000;
      coeffs_in_data_log_force[3418] <= 16'h0000;
      coeffs_in_data_log_force[3419] <= 16'h0000;
      coeffs_in_data_log_force[3420] <= 16'h0000;
      coeffs_in_data_log_force[3421] <= 16'h0000;
      coeffs_in_data_log_force[3422] <= 16'h0000;
      coeffs_in_data_log_force[3423] <= 16'h0000;
      coeffs_in_data_log_force[3424] <= 16'h0000;
      coeffs_in_data_log_force[3425] <= 16'h0000;
      coeffs_in_data_log_force[3426] <= 16'h0000;
      coeffs_in_data_log_force[3427] <= 16'h0000;
      coeffs_in_data_log_force[3428] <= 16'h0000;
      coeffs_in_data_log_force[3429] <= 16'h0000;
      coeffs_in_data_log_force[3430] <= 16'h0000;
      coeffs_in_data_log_force[3431] <= 16'h0000;
      coeffs_in_data_log_force[3432] <= 16'h0000;
      coeffs_in_data_log_force[3433] <= 16'h0000;
      coeffs_in_data_log_force[3434] <= 16'h0000;
      coeffs_in_data_log_force[3435] <= 16'h0000;
      coeffs_in_data_log_force[3436] <= 16'h0000;
      coeffs_in_data_log_force[3437] <= 16'h0000;
      coeffs_in_data_log_force[3438] <= 16'h0000;
      coeffs_in_data_log_force[3439] <= 16'h0000;
      coeffs_in_data_log_force[3440] <= 16'h0000;
      coeffs_in_data_log_force[3441] <= 16'h0000;
      coeffs_in_data_log_force[3442] <= 16'h0000;
      coeffs_in_data_log_force[3443] <= 16'h0000;
      coeffs_in_data_log_force[3444] <= 16'h0000;
      coeffs_in_data_log_force[3445] <= 16'h0000;
      coeffs_in_data_log_force[3446] <= 16'h0000;
      coeffs_in_data_log_force[3447] <= 16'h0000;
      coeffs_in_data_log_force[3448] <= 16'h0000;
      coeffs_in_data_log_force[3449] <= 16'h0000;
      coeffs_in_data_log_force[3450] <= 16'h0000;
      coeffs_in_data_log_force[3451] <= 16'h0000;
      coeffs_in_data_log_force[3452] <= 16'h0000;
      coeffs_in_data_log_force[3453] <= 16'h0000;
      coeffs_in_data_log_force[3454] <= 16'h0000;
      coeffs_in_data_log_force[3455] <= 16'h0000;
      coeffs_in_data_log_force[3456] <= 16'h0000;
      coeffs_in_data_log_force[3457] <= 16'h0000;
      coeffs_in_data_log_force[3458] <= 16'h0000;
      coeffs_in_data_log_force[3459] <= 16'h0000;
      coeffs_in_data_log_force[3460] <= 16'h0000;
      coeffs_in_data_log_force[3461] <= 16'h0000;
      coeffs_in_data_log_force[3462] <= 16'h0000;
      coeffs_in_data_log_force[3463] <= 16'h0000;
      coeffs_in_data_log_force[3464] <= 16'h0000;
      coeffs_in_data_log_force[3465] <= 16'h0000;
      coeffs_in_data_log_force[3466] <= 16'h0000;
      coeffs_in_data_log_force[3467] <= 16'h0000;
      coeffs_in_data_log_force[3468] <= 16'h0000;
      coeffs_in_data_log_force[3469] <= 16'h0000;
      coeffs_in_data_log_force[3470] <= 16'h0000;
      coeffs_in_data_log_force[3471] <= 16'h0000;
      coeffs_in_data_log_force[3472] <= 16'h0000;
      coeffs_in_data_log_force[3473] <= 16'h0000;
      coeffs_in_data_log_force[3474] <= 16'h0000;
      coeffs_in_data_log_force[3475] <= 16'h0000;
      coeffs_in_data_log_force[3476] <= 16'h0000;
      coeffs_in_data_log_force[3477] <= 16'h0000;
      coeffs_in_data_log_force[3478] <= 16'h0000;
      coeffs_in_data_log_force[3479] <= 16'h0000;
      coeffs_in_data_log_force[3480] <= 16'h0000;
      coeffs_in_data_log_force[3481] <= 16'h0000;
      coeffs_in_data_log_force[3482] <= 16'h0000;
      coeffs_in_data_log_force[3483] <= 16'h0000;
      coeffs_in_data_log_force[3484] <= 16'h0000;
      coeffs_in_data_log_force[3485] <= 16'h0000;
      coeffs_in_data_log_force[3486] <= 16'h0000;
      coeffs_in_data_log_force[3487] <= 16'h0000;
      coeffs_in_data_log_force[3488] <= 16'h0000;
      coeffs_in_data_log_force[3489] <= 16'h0000;
      coeffs_in_data_log_force[3490] <= 16'h0000;
      coeffs_in_data_log_force[3491] <= 16'h0000;
      coeffs_in_data_log_force[3492] <= 16'h0000;
      coeffs_in_data_log_force[3493] <= 16'h0000;
      coeffs_in_data_log_force[3494] <= 16'h0000;
      coeffs_in_data_log_force[3495] <= 16'h0000;
      coeffs_in_data_log_force[3496] <= 16'h0000;
      coeffs_in_data_log_force[3497] <= 16'h0000;
      coeffs_in_data_log_force[3498] <= 16'h0000;
      coeffs_in_data_log_force[3499] <= 16'h0000;
      coeffs_in_data_log_force[3500] <= 16'h0000;
      coeffs_in_data_log_force[3501] <= 16'h0000;
      coeffs_in_data_log_force[3502] <= 16'h0000;
      coeffs_in_data_log_force[3503] <= 16'h0000;
      coeffs_in_data_log_force[3504] <= 16'h0000;
      coeffs_in_data_log_force[3505] <= 16'h0000;
      coeffs_in_data_log_force[3506] <= 16'h0000;
      coeffs_in_data_log_force[3507] <= 16'h0000;
      coeffs_in_data_log_force[3508] <= 16'h0000;
      coeffs_in_data_log_force[3509] <= 16'h0000;
      coeffs_in_data_log_force[3510] <= 16'h0000;
      coeffs_in_data_log_force[3511] <= 16'h0000;
      coeffs_in_data_log_force[3512] <= 16'h0000;
      coeffs_in_data_log_force[3513] <= 16'h0000;
      coeffs_in_data_log_force[3514] <= 16'h0000;
      coeffs_in_data_log_force[3515] <= 16'h0000;
      coeffs_in_data_log_force[3516] <= 16'h0000;
      coeffs_in_data_log_force[3517] <= 16'h0000;
      coeffs_in_data_log_force[3518] <= 16'h0000;
      coeffs_in_data_log_force[3519] <= 16'h0000;
      coeffs_in_data_log_force[3520] <= 16'h0000;
      coeffs_in_data_log_force[3521] <= 16'h0000;
      coeffs_in_data_log_force[3522] <= 16'h0000;
      coeffs_in_data_log_force[3523] <= 16'h0000;
      coeffs_in_data_log_force[3524] <= 16'h0000;
      coeffs_in_data_log_force[3525] <= 16'h0000;
      coeffs_in_data_log_force[3526] <= 16'h0000;
      coeffs_in_data_log_force[3527] <= 16'h0000;
      coeffs_in_data_log_force[3528] <= 16'h0000;
      coeffs_in_data_log_force[3529] <= 16'h0000;
      coeffs_in_data_log_force[3530] <= 16'h0000;
      coeffs_in_data_log_force[3531] <= 16'h0000;
      coeffs_in_data_log_force[3532] <= 16'h0000;
      coeffs_in_data_log_force[3533] <= 16'h0000;
      coeffs_in_data_log_force[3534] <= 16'h0000;
      coeffs_in_data_log_force[3535] <= 16'h0000;
      coeffs_in_data_log_force[3536] <= 16'h0000;
      coeffs_in_data_log_force[3537] <= 16'h0000;
      coeffs_in_data_log_force[3538] <= 16'h0000;
      coeffs_in_data_log_force[3539] <= 16'h0000;
      coeffs_in_data_log_force[3540] <= 16'h0000;
      coeffs_in_data_log_force[3541] <= 16'h0000;
      coeffs_in_data_log_force[3542] <= 16'h0000;
      coeffs_in_data_log_force[3543] <= 16'h0000;
      coeffs_in_data_log_force[3544] <= 16'h0000;
      coeffs_in_data_log_force[3545] <= 16'h0000;
      coeffs_in_data_log_force[3546] <= 16'h0000;
      coeffs_in_data_log_force[3547] <= 16'h0000;
      coeffs_in_data_log_force[3548] <= 16'h0000;
      coeffs_in_data_log_force[3549] <= 16'h0000;
      coeffs_in_data_log_force[3550] <= 16'h0000;
      coeffs_in_data_log_force[3551] <= 16'h0000;
      coeffs_in_data_log_force[3552] <= 16'h0000;
      coeffs_in_data_log_force[3553] <= 16'h0000;
      coeffs_in_data_log_force[3554] <= 16'h0000;
      coeffs_in_data_log_force[3555] <= 16'h0000;
      coeffs_in_data_log_force[3556] <= 16'h0000;
      coeffs_in_data_log_force[3557] <= 16'h0000;
      coeffs_in_data_log_force[3558] <= 16'h0000;
      coeffs_in_data_log_force[3559] <= 16'h0000;
      coeffs_in_data_log_force[3560] <= 16'h0000;
      coeffs_in_data_log_force[3561] <= 16'h0000;
      coeffs_in_data_log_force[3562] <= 16'h0000;
      coeffs_in_data_log_force[3563] <= 16'h0000;
      coeffs_in_data_log_force[3564] <= 16'h0000;
      coeffs_in_data_log_force[3565] <= 16'h0000;
      coeffs_in_data_log_force[3566] <= 16'h0000;
      coeffs_in_data_log_force[3567] <= 16'h0000;
      coeffs_in_data_log_force[3568] <= 16'h0000;
      coeffs_in_data_log_force[3569] <= 16'h0000;
      coeffs_in_data_log_force[3570] <= 16'h0000;
      coeffs_in_data_log_force[3571] <= 16'h0000;
      coeffs_in_data_log_force[3572] <= 16'h0000;
      coeffs_in_data_log_force[3573] <= 16'h0000;
      coeffs_in_data_log_force[3574] <= 16'h0000;
      coeffs_in_data_log_force[3575] <= 16'h0000;
      coeffs_in_data_log_force[3576] <= 16'h0000;
      coeffs_in_data_log_force[3577] <= 16'h0000;
      coeffs_in_data_log_force[3578] <= 16'h0000;
      coeffs_in_data_log_force[3579] <= 16'h0000;
      coeffs_in_data_log_force[3580] <= 16'h0000;
      coeffs_in_data_log_force[3581] <= 16'h0000;
      coeffs_in_data_log_force[3582] <= 16'h0000;
      coeffs_in_data_log_force[3583] <= 16'h0000;
      coeffs_in_data_log_force[3584] <= 16'h0000;
      coeffs_in_data_log_force[3585] <= 16'h0000;
      coeffs_in_data_log_force[3586] <= 16'h0000;
      coeffs_in_data_log_force[3587] <= 16'h0000;
      coeffs_in_data_log_force[3588] <= 16'h0000;
      coeffs_in_data_log_force[3589] <= 16'h0000;
      coeffs_in_data_log_force[3590] <= 16'h0000;
      coeffs_in_data_log_force[3591] <= 16'h0000;
      coeffs_in_data_log_force[3592] <= 16'h0000;
      coeffs_in_data_log_force[3593] <= 16'h0000;
      coeffs_in_data_log_force[3594] <= 16'h0000;
      coeffs_in_data_log_force[3595] <= 16'h0000;
      coeffs_in_data_log_force[3596] <= 16'h0000;
      coeffs_in_data_log_force[3597] <= 16'h0000;
      coeffs_in_data_log_force[3598] <= 16'h0000;
      coeffs_in_data_log_force[3599] <= 16'h0000;
      coeffs_in_data_log_force[3600] <= 16'h0000;
      coeffs_in_data_log_force[3601] <= 16'h0000;
      coeffs_in_data_log_force[3602] <= 16'h0000;
      coeffs_in_data_log_force[3603] <= 16'h0000;
      coeffs_in_data_log_force[3604] <= 16'h0000;
      coeffs_in_data_log_force[3605] <= 16'h0000;
      coeffs_in_data_log_force[3606] <= 16'h0000;
      coeffs_in_data_log_force[3607] <= 16'h0000;
      coeffs_in_data_log_force[3608] <= 16'h0000;
      coeffs_in_data_log_force[3609] <= 16'h0000;
      coeffs_in_data_log_force[3610] <= 16'h0000;
      coeffs_in_data_log_force[3611] <= 16'h0000;
      coeffs_in_data_log_force[3612] <= 16'h0000;
      coeffs_in_data_log_force[3613] <= 16'h0000;
      coeffs_in_data_log_force[3614] <= 16'h0000;
      coeffs_in_data_log_force[3615] <= 16'h0000;
      coeffs_in_data_log_force[3616] <= 16'h0000;
      coeffs_in_data_log_force[3617] <= 16'h0000;
      coeffs_in_data_log_force[3618] <= 16'h0000;
      coeffs_in_data_log_force[3619] <= 16'h0000;
      coeffs_in_data_log_force[3620] <= 16'h0000;
      coeffs_in_data_log_force[3621] <= 16'h0000;
      coeffs_in_data_log_force[3622] <= 16'h0000;
      coeffs_in_data_log_force[3623] <= 16'h0000;
      coeffs_in_data_log_force[3624] <= 16'h0000;
      coeffs_in_data_log_force[3625] <= 16'h0000;
      coeffs_in_data_log_force[3626] <= 16'h0000;
      coeffs_in_data_log_force[3627] <= 16'h0000;
      coeffs_in_data_log_force[3628] <= 16'h0000;
      coeffs_in_data_log_force[3629] <= 16'h0000;
      coeffs_in_data_log_force[3630] <= 16'h0000;
      coeffs_in_data_log_force[3631] <= 16'h0000;
      coeffs_in_data_log_force[3632] <= 16'h0000;
      coeffs_in_data_log_force[3633] <= 16'h0000;
      coeffs_in_data_log_force[3634] <= 16'h0000;
      coeffs_in_data_log_force[3635] <= 16'h0000;
      coeffs_in_data_log_force[3636] <= 16'h0000;
      coeffs_in_data_log_force[3637] <= 16'h0000;
      coeffs_in_data_log_force[3638] <= 16'h0000;
      coeffs_in_data_log_force[3639] <= 16'h0000;
      coeffs_in_data_log_force[3640] <= 16'h0000;
      coeffs_in_data_log_force[3641] <= 16'h0000;
      coeffs_in_data_log_force[3642] <= 16'h0000;
      coeffs_in_data_log_force[3643] <= 16'h0000;
      coeffs_in_data_log_force[3644] <= 16'h0000;
      coeffs_in_data_log_force[3645] <= 16'h0000;
      coeffs_in_data_log_force[3646] <= 16'h0000;
      coeffs_in_data_log_force[3647] <= 16'h0000;
      coeffs_in_data_log_force[3648] <= 16'h0000;
      coeffs_in_data_log_force[3649] <= 16'h0000;
      coeffs_in_data_log_force[3650] <= 16'h0000;
      coeffs_in_data_log_force[3651] <= 16'h0000;
      coeffs_in_data_log_force[3652] <= 16'h0000;
      coeffs_in_data_log_force[3653] <= 16'h0000;
      coeffs_in_data_log_force[3654] <= 16'h0000;
      coeffs_in_data_log_force[3655] <= 16'h0000;
      coeffs_in_data_log_force[3656] <= 16'h0000;
      coeffs_in_data_log_force[3657] <= 16'h0000;
      coeffs_in_data_log_force[3658] <= 16'h0000;
      coeffs_in_data_log_force[3659] <= 16'h0000;
      coeffs_in_data_log_force[3660] <= 16'h0000;
      coeffs_in_data_log_force[3661] <= 16'h0000;
      coeffs_in_data_log_force[3662] <= 16'h0000;
      coeffs_in_data_log_force[3663] <= 16'h0000;
      coeffs_in_data_log_force[3664] <= 16'h0000;
      coeffs_in_data_log_force[3665] <= 16'h0000;
      coeffs_in_data_log_force[3666] <= 16'h0000;
      coeffs_in_data_log_force[3667] <= 16'h0000;
      coeffs_in_data_log_force[3668] <= 16'h0000;
      coeffs_in_data_log_force[3669] <= 16'h0000;
      coeffs_in_data_log_force[3670] <= 16'h0000;
      coeffs_in_data_log_force[3671] <= 16'h0000;
      coeffs_in_data_log_force[3672] <= 16'h0000;
      coeffs_in_data_log_force[3673] <= 16'h0000;
      coeffs_in_data_log_force[3674] <= 16'h0000;
      coeffs_in_data_log_force[3675] <= 16'h0000;
      coeffs_in_data_log_force[3676] <= 16'h0000;
      coeffs_in_data_log_force[3677] <= 16'h0000;
      coeffs_in_data_log_force[3678] <= 16'h0000;
      coeffs_in_data_log_force[3679] <= 16'h0000;
      coeffs_in_data_log_force[3680] <= 16'h0000;
      coeffs_in_data_log_force[3681] <= 16'h0000;
      coeffs_in_data_log_force[3682] <= 16'h0000;
      coeffs_in_data_log_force[3683] <= 16'h0000;
      coeffs_in_data_log_force[3684] <= 16'h0000;
      coeffs_in_data_log_force[3685] <= 16'h0000;
      coeffs_in_data_log_force[3686] <= 16'h0000;
      coeffs_in_data_log_force[3687] <= 16'h0000;
      coeffs_in_data_log_force[3688] <= 16'h0000;
      coeffs_in_data_log_force[3689] <= 16'h0000;
      coeffs_in_data_log_force[3690] <= 16'h0000;
      coeffs_in_data_log_force[3691] <= 16'h0000;
      coeffs_in_data_log_force[3692] <= 16'h0000;
      coeffs_in_data_log_force[3693] <= 16'h0000;
      coeffs_in_data_log_force[3694] <= 16'h0000;
      coeffs_in_data_log_force[3695] <= 16'h0000;
      coeffs_in_data_log_force[3696] <= 16'h0000;
      coeffs_in_data_log_force[3697] <= 16'h0000;
      coeffs_in_data_log_force[3698] <= 16'h0000;
      coeffs_in_data_log_force[3699] <= 16'h0000;
      coeffs_in_data_log_force[3700] <= 16'h0000;
      coeffs_in_data_log_force[3701] <= 16'h0000;
      coeffs_in_data_log_force[3702] <= 16'h0000;
      coeffs_in_data_log_force[3703] <= 16'h0000;
      coeffs_in_data_log_force[3704] <= 16'h0000;
      coeffs_in_data_log_force[3705] <= 16'h0000;
      coeffs_in_data_log_force[3706] <= 16'h0000;
      coeffs_in_data_log_force[3707] <= 16'h0000;
      coeffs_in_data_log_force[3708] <= 16'h0000;
      coeffs_in_data_log_force[3709] <= 16'h0000;
      coeffs_in_data_log_force[3710] <= 16'h0000;
      coeffs_in_data_log_force[3711] <= 16'h0000;
      coeffs_in_data_log_force[3712] <= 16'h0000;
      coeffs_in_data_log_force[3713] <= 16'h0000;
      coeffs_in_data_log_force[3714] <= 16'h0000;
      coeffs_in_data_log_force[3715] <= 16'h0000;
      coeffs_in_data_log_force[3716] <= 16'h0000;
      coeffs_in_data_log_force[3717] <= 16'h0000;
      coeffs_in_data_log_force[3718] <= 16'h0000;
      coeffs_in_data_log_force[3719] <= 16'h0000;
      coeffs_in_data_log_force[3720] <= 16'h0000;
      coeffs_in_data_log_force[3721] <= 16'h0000;
      coeffs_in_data_log_force[3722] <= 16'h0000;
      coeffs_in_data_log_force[3723] <= 16'h0000;
      coeffs_in_data_log_force[3724] <= 16'h0000;
      coeffs_in_data_log_force[3725] <= 16'h0000;
      coeffs_in_data_log_force[3726] <= 16'h0000;
      coeffs_in_data_log_force[3727] <= 16'h0000;
      coeffs_in_data_log_force[3728] <= 16'h0000;
      coeffs_in_data_log_force[3729] <= 16'h0000;
      coeffs_in_data_log_force[3730] <= 16'h0000;
      coeffs_in_data_log_force[3731] <= 16'h0000;
      coeffs_in_data_log_force[3732] <= 16'h0000;
      coeffs_in_data_log_force[3733] <= 16'h0000;
      coeffs_in_data_log_force[3734] <= 16'h0000;
      coeffs_in_data_log_force[3735] <= 16'h0000;
      coeffs_in_data_log_force[3736] <= 16'h0000;
      coeffs_in_data_log_force[3737] <= 16'h0000;
      coeffs_in_data_log_force[3738] <= 16'h0000;
      coeffs_in_data_log_force[3739] <= 16'h0000;
      coeffs_in_data_log_force[3740] <= 16'h0000;
      coeffs_in_data_log_force[3741] <= 16'h0000;
      coeffs_in_data_log_force[3742] <= 16'h0000;
      coeffs_in_data_log_force[3743] <= 16'h0000;
      coeffs_in_data_log_force[3744] <= 16'h0000;
      coeffs_in_data_log_force[3745] <= 16'h0000;
      coeffs_in_data_log_force[3746] <= 16'h0000;
      coeffs_in_data_log_force[3747] <= 16'h0000;
      coeffs_in_data_log_force[3748] <= 16'h0000;
      coeffs_in_data_log_force[3749] <= 16'h0000;
      coeffs_in_data_log_force[3750] <= 16'h0000;
      coeffs_in_data_log_force[3751] <= 16'h0000;
      coeffs_in_data_log_force[3752] <= 16'h0000;
      coeffs_in_data_log_force[3753] <= 16'h0000;
      coeffs_in_data_log_force[3754] <= 16'h0000;
      coeffs_in_data_log_force[3755] <= 16'h0000;
      coeffs_in_data_log_force[3756] <= 16'h0000;
      coeffs_in_data_log_force[3757] <= 16'h0000;
      coeffs_in_data_log_force[3758] <= 16'h0000;
      coeffs_in_data_log_force[3759] <= 16'h0000;
      coeffs_in_data_log_force[3760] <= 16'h0000;
      coeffs_in_data_log_force[3761] <= 16'h0000;
      coeffs_in_data_log_force[3762] <= 16'h0000;
      coeffs_in_data_log_force[3763] <= 16'h0000;
      coeffs_in_data_log_force[3764] <= 16'h0000;
      coeffs_in_data_log_force[3765] <= 16'h0000;
      coeffs_in_data_log_force[3766] <= 16'h0000;
      coeffs_in_data_log_force[3767] <= 16'h0000;
      coeffs_in_data_log_force[3768] <= 16'h0000;
      coeffs_in_data_log_force[3769] <= 16'h0000;
      coeffs_in_data_log_force[3770] <= 16'h0000;
      coeffs_in_data_log_force[3771] <= 16'h0000;
      coeffs_in_data_log_force[3772] <= 16'h0000;
      coeffs_in_data_log_force[3773] <= 16'h0000;
      coeffs_in_data_log_force[3774] <= 16'h0000;
      coeffs_in_data_log_force[3775] <= 16'h0000;
      coeffs_in_data_log_force[3776] <= 16'h0000;
      coeffs_in_data_log_force[3777] <= 16'h0000;
      coeffs_in_data_log_force[3778] <= 16'h0000;
      coeffs_in_data_log_force[3779] <= 16'h0000;
      coeffs_in_data_log_force[3780] <= 16'h0000;
      coeffs_in_data_log_force[3781] <= 16'h0000;
      coeffs_in_data_log_force[3782] <= 16'h0000;
      coeffs_in_data_log_force[3783] <= 16'h0000;
      coeffs_in_data_log_force[3784] <= 16'h0000;
      coeffs_in_data_log_force[3785] <= 16'h0000;
      coeffs_in_data_log_force[3786] <= 16'h0000;
      coeffs_in_data_log_force[3787] <= 16'h0000;
      coeffs_in_data_log_force[3788] <= 16'h0000;
      coeffs_in_data_log_force[3789] <= 16'h0000;
      coeffs_in_data_log_force[3790] <= 16'h0000;
      coeffs_in_data_log_force[3791] <= 16'h0000;
      coeffs_in_data_log_force[3792] <= 16'h0000;
      coeffs_in_data_log_force[3793] <= 16'h0000;
      coeffs_in_data_log_force[3794] <= 16'h0000;
      coeffs_in_data_log_force[3795] <= 16'h0000;
      coeffs_in_data_log_force[3796] <= 16'h0000;
      coeffs_in_data_log_force[3797] <= 16'h0000;
      coeffs_in_data_log_force[3798] <= 16'h0000;
      coeffs_in_data_log_force[3799] <= 16'h0000;
      coeffs_in_data_log_force[3800] <= 16'h0000;
      coeffs_in_data_log_force[3801] <= 16'h0000;
      coeffs_in_data_log_force[3802] <= 16'h0000;
      coeffs_in_data_log_force[3803] <= 16'h0000;
      coeffs_in_data_log_force[3804] <= 16'h0000;
      coeffs_in_data_log_force[3805] <= 16'h0000;
      coeffs_in_data_log_force[3806] <= 16'h0000;
      coeffs_in_data_log_force[3807] <= 16'h0000;
      coeffs_in_data_log_force[3808] <= 16'h0000;
      coeffs_in_data_log_force[3809] <= 16'h0000;
      coeffs_in_data_log_force[3810] <= 16'h0000;
      coeffs_in_data_log_force[3811] <= 16'h0000;
      coeffs_in_data_log_force[3812] <= 16'h0000;
      coeffs_in_data_log_force[3813] <= 16'h0000;
      coeffs_in_data_log_force[3814] <= 16'h0000;
      coeffs_in_data_log_force[3815] <= 16'h0000;
      coeffs_in_data_log_force[3816] <= 16'h0000;
      coeffs_in_data_log_force[3817] <= 16'h0000;
      coeffs_in_data_log_force[3818] <= 16'h0000;
      coeffs_in_data_log_force[3819] <= 16'h0000;
      coeffs_in_data_log_force[3820] <= 16'h0000;
      coeffs_in_data_log_force[3821] <= 16'h0000;
      coeffs_in_data_log_force[3822] <= 16'h0000;
      coeffs_in_data_log_force[3823] <= 16'h0000;
      coeffs_in_data_log_force[3824] <= 16'h0000;
      coeffs_in_data_log_force[3825] <= 16'h0000;
      coeffs_in_data_log_force[3826] <= 16'h0000;
      coeffs_in_data_log_force[3827] <= 16'h0000;
      coeffs_in_data_log_force[3828] <= 16'h0000;
      coeffs_in_data_log_force[3829] <= 16'h0000;
      coeffs_in_data_log_force[3830] <= 16'h0000;
      coeffs_in_data_log_force[3831] <= 16'h0000;
      coeffs_in_data_log_force[3832] <= 16'h0000;
      coeffs_in_data_log_force[3833] <= 16'h0000;
      coeffs_in_data_log_force[3834] <= 16'h0000;
      coeffs_in_data_log_force[3835] <= 16'h0000;
      coeffs_in_data_log_force[3836] <= 16'h0000;
      coeffs_in_data_log_force[3837] <= 16'h0000;
      coeffs_in_data_log_force[3838] <= 16'h0000;
      coeffs_in_data_log_force[3839] <= 16'h0000;
      coeffs_in_data_log_force[3840] <= 16'h0000;
      coeffs_in_data_log_force[3841] <= 16'h0000;
      coeffs_in_data_log_force[3842] <= 16'h0000;
      coeffs_in_data_log_force[3843] <= 16'h0000;
      coeffs_in_data_log_force[3844] <= 16'h0000;
      coeffs_in_data_log_force[3845] <= 16'h0000;
      coeffs_in_data_log_force[3846] <= 16'h0000;
      coeffs_in_data_log_force[3847] <= 16'h0000;
      coeffs_in_data_log_force[3848] <= 16'h0000;
      coeffs_in_data_log_force[3849] <= 16'h0000;
      coeffs_in_data_log_force[3850] <= 16'h0000;
      coeffs_in_data_log_force[3851] <= 16'h0000;
      coeffs_in_data_log_force[3852] <= 16'h0000;
      coeffs_in_data_log_force[3853] <= 16'h0000;
      coeffs_in_data_log_force[3854] <= 16'h0000;
      coeffs_in_data_log_force[3855] <= 16'h0000;
      coeffs_in_data_log_force[3856] <= 16'h0000;
      coeffs_in_data_log_force[3857] <= 16'h0000;
      coeffs_in_data_log_force[3858] <= 16'h0000;
      coeffs_in_data_log_force[3859] <= 16'h0000;
      coeffs_in_data_log_force[3860] <= 16'h0000;
      coeffs_in_data_log_force[3861] <= 16'h0000;
      coeffs_in_data_log_force[3862] <= 16'h0000;
      coeffs_in_data_log_force[3863] <= 16'h0000;
      coeffs_in_data_log_force[3864] <= 16'h0000;
      coeffs_in_data_log_force[3865] <= 16'h0000;
      coeffs_in_data_log_force[3866] <= 16'h0000;
      coeffs_in_data_log_force[3867] <= 16'h0000;
      coeffs_in_data_log_force[3868] <= 16'h0000;
      coeffs_in_data_log_force[3869] <= 16'h0000;
      coeffs_in_data_log_force[3870] <= 16'h0000;
      coeffs_in_data_log_force[3871] <= 16'h0000;
      coeffs_in_data_log_force[3872] <= 16'h0000;
      coeffs_in_data_log_force[3873] <= 16'h0000;
      coeffs_in_data_log_force[3874] <= 16'h0000;
      coeffs_in_data_log_force[3875] <= 16'h0000;
      coeffs_in_data_log_force[3876] <= 16'h0000;
      coeffs_in_data_log_force[3877] <= 16'h0000;
      coeffs_in_data_log_force[3878] <= 16'h0000;
      coeffs_in_data_log_force[3879] <= 16'h0000;
      coeffs_in_data_log_force[3880] <= 16'h0000;
      coeffs_in_data_log_force[3881] <= 16'h0000;
      coeffs_in_data_log_force[3882] <= 16'h0000;
      coeffs_in_data_log_force[3883] <= 16'h0000;
      coeffs_in_data_log_force[3884] <= 16'h0000;
      coeffs_in_data_log_force[3885] <= 16'h0000;
      coeffs_in_data_log_force[3886] <= 16'h0000;
      coeffs_in_data_log_force[3887] <= 16'h0000;
      coeffs_in_data_log_force[3888] <= 16'h0000;
      coeffs_in_data_log_force[3889] <= 16'h0000;
      coeffs_in_data_log_force[3890] <= 16'h0000;
      coeffs_in_data_log_force[3891] <= 16'h0000;
      coeffs_in_data_log_force[3892] <= 16'h0000;
      coeffs_in_data_log_force[3893] <= 16'h0000;
      coeffs_in_data_log_force[3894] <= 16'h0000;
      coeffs_in_data_log_force[3895] <= 16'h0000;
      coeffs_in_data_log_force[3896] <= 16'h0000;
      coeffs_in_data_log_force[3897] <= 16'h0000;
      coeffs_in_data_log_force[3898] <= 16'h0000;
      coeffs_in_data_log_force[3899] <= 16'h0000;
      coeffs_in_data_log_force[3900] <= 16'h0000;
      coeffs_in_data_log_force[3901] <= 16'h0000;
      coeffs_in_data_log_force[3902] <= 16'h0000;
      coeffs_in_data_log_force[3903] <= 16'h0000;
      coeffs_in_data_log_force[3904] <= 16'h0000;
      coeffs_in_data_log_force[3905] <= 16'h0000;
      coeffs_in_data_log_force[3906] <= 16'h0000;
      coeffs_in_data_log_force[3907] <= 16'h0000;
      coeffs_in_data_log_force[3908] <= 16'h0000;
      coeffs_in_data_log_force[3909] <= 16'h0000;
      coeffs_in_data_log_force[3910] <= 16'h0000;
      coeffs_in_data_log_force[3911] <= 16'h0000;
      coeffs_in_data_log_force[3912] <= 16'h0000;
      coeffs_in_data_log_force[3913] <= 16'h0000;
      coeffs_in_data_log_force[3914] <= 16'h0000;
      coeffs_in_data_log_force[3915] <= 16'h0000;
      coeffs_in_data_log_force[3916] <= 16'h0000;
      coeffs_in_data_log_force[3917] <= 16'h0000;
      coeffs_in_data_log_force[3918] <= 16'h0000;
      coeffs_in_data_log_force[3919] <= 16'h0000;
      coeffs_in_data_log_force[3920] <= 16'h0000;
      coeffs_in_data_log_force[3921] <= 16'h0000;
      coeffs_in_data_log_force[3922] <= 16'h0000;
      coeffs_in_data_log_force[3923] <= 16'h0000;
      coeffs_in_data_log_force[3924] <= 16'h0000;
      coeffs_in_data_log_force[3925] <= 16'h0000;
      coeffs_in_data_log_force[3926] <= 16'h0000;
      coeffs_in_data_log_force[3927] <= 16'h0000;
      coeffs_in_data_log_force[3928] <= 16'h0000;
      coeffs_in_data_log_force[3929] <= 16'h0000;
      coeffs_in_data_log_force[3930] <= 16'h0000;
      coeffs_in_data_log_force[3931] <= 16'h0000;
      coeffs_in_data_log_force[3932] <= 16'h0000;
      coeffs_in_data_log_force[3933] <= 16'h0000;
      coeffs_in_data_log_force[3934] <= 16'h0000;
      coeffs_in_data_log_force[3935] <= 16'h0000;
      coeffs_in_data_log_force[3936] <= 16'h0000;
      coeffs_in_data_log_force[3937] <= 16'h0000;
      coeffs_in_data_log_force[3938] <= 16'h0000;
      coeffs_in_data_log_force[3939] <= 16'h0000;
      coeffs_in_data_log_force[3940] <= 16'h0000;
      coeffs_in_data_log_force[3941] <= 16'h0000;
      coeffs_in_data_log_force[3942] <= 16'h0000;
      coeffs_in_data_log_force[3943] <= 16'h0000;
      coeffs_in_data_log_force[3944] <= 16'h0000;
      coeffs_in_data_log_force[3945] <= 16'h0000;
      coeffs_in_data_log_force[3946] <= 16'h0000;
      coeffs_in_data_log_force[3947] <= 16'h0000;
      coeffs_in_data_log_force[3948] <= 16'h0000;
      coeffs_in_data_log_force[3949] <= 16'h0000;
      coeffs_in_data_log_force[3950] <= 16'h0000;
      coeffs_in_data_log_force[3951] <= 16'h0000;
      coeffs_in_data_log_force[3952] <= 16'h0000;
      coeffs_in_data_log_force[3953] <= 16'h0000;
      coeffs_in_data_log_force[3954] <= 16'h0000;
      coeffs_in_data_log_force[3955] <= 16'h0000;
      coeffs_in_data_log_force[3956] <= 16'h0000;
      coeffs_in_data_log_force[3957] <= 16'h0000;
      coeffs_in_data_log_force[3958] <= 16'h0000;
      coeffs_in_data_log_force[3959] <= 16'h0000;
      coeffs_in_data_log_force[3960] <= 16'h0000;
      coeffs_in_data_log_force[3961] <= 16'h0000;
      coeffs_in_data_log_force[3962] <= 16'h0000;
      coeffs_in_data_log_force[3963] <= 16'h0000;
      coeffs_in_data_log_force[3964] <= 16'h0000;
      coeffs_in_data_log_force[3965] <= 16'h0000;
      coeffs_in_data_log_force[3966] <= 16'h0000;
      coeffs_in_data_log_force[3967] <= 16'h0000;
      coeffs_in_data_log_force[3968] <= 16'h0000;
      coeffs_in_data_log_force[3969] <= 16'h0000;
      coeffs_in_data_log_force[3970] <= 16'h0000;
      coeffs_in_data_log_force[3971] <= 16'h0000;
      coeffs_in_data_log_force[3972] <= 16'h0000;
      coeffs_in_data_log_force[3973] <= 16'h0000;
      coeffs_in_data_log_force[3974] <= 16'h0000;
      coeffs_in_data_log_force[3975] <= 16'h0000;
      coeffs_in_data_log_force[3976] <= 16'h0000;
      coeffs_in_data_log_force[3977] <= 16'h0000;
      coeffs_in_data_log_force[3978] <= 16'h0000;
      coeffs_in_data_log_force[3979] <= 16'h0000;
      coeffs_in_data_log_force[3980] <= 16'h0000;
      coeffs_in_data_log_force[3981] <= 16'h0000;
      coeffs_in_data_log_force[3982] <= 16'h0000;
      coeffs_in_data_log_force[3983] <= 16'h0000;
      coeffs_in_data_log_force[3984] <= 16'h0000;
      coeffs_in_data_log_force[3985] <= 16'h0000;
      coeffs_in_data_log_force[3986] <= 16'h0000;
      coeffs_in_data_log_force[3987] <= 16'h0000;
      coeffs_in_data_log_force[3988] <= 16'h0000;
      coeffs_in_data_log_force[3989] <= 16'h0000;
      coeffs_in_data_log_force[3990] <= 16'h0000;
      coeffs_in_data_log_force[3991] <= 16'h0000;
      coeffs_in_data_log_force[3992] <= 16'h0000;
      coeffs_in_data_log_force[3993] <= 16'h0000;
      coeffs_in_data_log_force[3994] <= 16'h0000;
      coeffs_in_data_log_force[3995] <= 16'h0000;
      coeffs_in_data_log_force[3996] <= 16'h0000;
      coeffs_in_data_log_force[3997] <= 16'h0000;
      coeffs_in_data_log_force[3998] <= 16'h0000;
      coeffs_in_data_log_force[3999] <= 16'h0000;
      coeffs_in_data_log_force[4000] <= 16'h0000;
      coeffs_in_data_log_force[4001] <= 16'h0000;
      coeffs_in_data_log_force[4002] <= 16'h0000;
      coeffs_in_data_log_force[4003] <= 16'h0000;
      coeffs_in_data_log_force[4004] <= 16'h0000;
      coeffs_in_data_log_force[4005] <= 16'h0000;
      coeffs_in_data_log_force[4006] <= 16'h0000;
      coeffs_in_data_log_force[4007] <= 16'h0000;
      coeffs_in_data_log_force[4008] <= 16'h0000;
      coeffs_in_data_log_force[4009] <= 16'h0000;
      coeffs_in_data_log_force[4010] <= 16'h0000;
      coeffs_in_data_log_force[4011] <= 16'h0000;
      coeffs_in_data_log_force[4012] <= 16'h0000;
      coeffs_in_data_log_force[4013] <= 16'h0000;
      coeffs_in_data_log_force[4014] <= 16'h0000;
      coeffs_in_data_log_force[4015] <= 16'h0000;
      coeffs_in_data_log_force[4016] <= 16'h0000;
      coeffs_in_data_log_force[4017] <= 16'h0000;
      coeffs_in_data_log_force[4018] <= 16'h0000;
      coeffs_in_data_log_force[4019] <= 16'h0000;
      coeffs_in_data_log_force[4020] <= 16'h0000;
      coeffs_in_data_log_force[4021] <= 16'h0000;
      coeffs_in_data_log_force[4022] <= 16'h0000;
      coeffs_in_data_log_force[4023] <= 16'h0000;
      coeffs_in_data_log_force[4024] <= 16'h0000;
      coeffs_in_data_log_force[4025] <= 16'h0000;
      coeffs_in_data_log_force[4026] <= 16'h0000;
      coeffs_in_data_log_force[4027] <= 16'h0000;
      coeffs_in_data_log_force[4028] <= 16'h0000;
      coeffs_in_data_log_force[4029] <= 16'h0000;
      coeffs_in_data_log_force[4030] <= 16'h0000;
      coeffs_in_data_log_force[4031] <= 16'h0000;
      coeffs_in_data_log_force[4032] <= 16'h0000;
      coeffs_in_data_log_force[4033] <= 16'h0000;
      coeffs_in_data_log_force[4034] <= 16'h0000;
      coeffs_in_data_log_force[4035] <= 16'h0000;
      coeffs_in_data_log_force[4036] <= 16'h0000;
      coeffs_in_data_log_force[4037] <= 16'h0000;
      coeffs_in_data_log_force[4038] <= 16'h0000;
      coeffs_in_data_log_force[4039] <= 16'h0000;
      coeffs_in_data_log_force[4040] <= 16'h0000;
      coeffs_in_data_log_force[4041] <= 16'h0000;
      coeffs_in_data_log_force[4042] <= 16'h0000;
      coeffs_in_data_log_force[4043] <= 16'h0000;
      coeffs_in_data_log_force[4044] <= 16'h0000;
      coeffs_in_data_log_force[4045] <= 16'h0000;
      coeffs_in_data_log_force[4046] <= 16'h0000;
      coeffs_in_data_log_force[4047] <= 16'h0000;
      coeffs_in_data_log_force[4048] <= 16'h0000;
      coeffs_in_data_log_force[4049] <= 16'h0000;
      coeffs_in_data_log_force[4050] <= 16'h0000;
      coeffs_in_data_log_force[4051] <= 16'h0000;
      coeffs_in_data_log_force[4052] <= 16'h0000;
      coeffs_in_data_log_force[4053] <= 16'h0000;
      coeffs_in_data_log_force[4054] <= 16'h0000;
      coeffs_in_data_log_force[4055] <= 16'h0000;
      coeffs_in_data_log_force[4056] <= 16'h0000;
      coeffs_in_data_log_force[4057] <= 16'h0000;
      coeffs_in_data_log_force[4058] <= 16'h0000;
      coeffs_in_data_log_force[4059] <= 16'h0000;
      coeffs_in_data_log_force[4060] <= 16'h0000;
      coeffs_in_data_log_force[4061] <= 16'h0000;
      coeffs_in_data_log_force[4062] <= 16'h0000;
      coeffs_in_data_log_force[4063] <= 16'h0000;
      coeffs_in_data_log_force[4064] <= 16'h0000;
      coeffs_in_data_log_force[4065] <= 16'h0000;
      coeffs_in_data_log_force[4066] <= 16'h0000;
      coeffs_in_data_log_force[4067] <= 16'h0000;
      coeffs_in_data_log_force[4068] <= 16'h0000;
      coeffs_in_data_log_force[4069] <= 16'h0000;
      coeffs_in_data_log_force[4070] <= 16'h0000;
      coeffs_in_data_log_force[4071] <= 16'h0000;
      coeffs_in_data_log_force[4072] <= 16'h0000;
      coeffs_in_data_log_force[4073] <= 16'h0000;
      coeffs_in_data_log_force[4074] <= 16'h0000;
      coeffs_in_data_log_force[4075] <= 16'h0000;
      coeffs_in_data_log_force[4076] <= 16'h0000;
      coeffs_in_data_log_force[4077] <= 16'h0000;
      coeffs_in_data_log_force[4078] <= 16'h0000;
      coeffs_in_data_log_force[4079] <= 16'h0000;
      coeffs_in_data_log_force[4080] <= 16'h0000;
      coeffs_in_data_log_force[4081] <= 16'h0000;
      coeffs_in_data_log_force[4082] <= 16'h0000;
      coeffs_in_data_log_force[4083] <= 16'h0000;
      coeffs_in_data_log_force[4084] <= 16'h0000;
      coeffs_in_data_log_force[4085] <= 16'h0000;
      coeffs_in_data_log_force[4086] <= 16'h0000;
      coeffs_in_data_log_force[4087] <= 16'h0000;
      coeffs_in_data_log_force[4088] <= 16'h0000;
      coeffs_in_data_log_force[4089] <= 16'h0000;
      coeffs_in_data_log_force[4090] <= 16'h0000;
      coeffs_in_data_log_force[4091] <= 16'h0000;
      coeffs_in_data_log_force[4092] <= 16'h0000;
      coeffs_in_data_log_force[4093] <= 16'h0000;
      coeffs_in_data_log_force[4094] <= 16'h0000;
      coeffs_in_data_log_force[4095] <= 16'h0000;
      coeffs_in_data_log_force[4096] <= 16'h0000;
      coeffs_in_data_log_force[4097] <= 16'h0000;
      coeffs_in_data_log_force[4098] <= 16'h0000;
      coeffs_in_data_log_force[4099] <= 16'h0000;
      coeffs_in_data_log_force[4100] <= 16'h0000;
      coeffs_in_data_log_force[4101] <= 16'h0000;
      coeffs_in_data_log_force[4102] <= 16'h0000;
      coeffs_in_data_log_force[4103] <= 16'h0000;
      coeffs_in_data_log_force[4104] <= 16'h0000;
      coeffs_in_data_log_force[4105] <= 16'h0000;
      coeffs_in_data_log_force[4106] <= 16'h0000;
      coeffs_in_data_log_force[4107] <= 16'h0000;
      coeffs_in_data_log_force[4108] <= 16'h0000;
      coeffs_in_data_log_force[4109] <= 16'h0000;
      coeffs_in_data_log_force[4110] <= 16'h0000;
      coeffs_in_data_log_force[4111] <= 16'h0000;
      coeffs_in_data_log_force[4112] <= 16'h0000;
      coeffs_in_data_log_force[4113] <= 16'h0000;
      coeffs_in_data_log_force[4114] <= 16'h0000;
      coeffs_in_data_log_force[4115] <= 16'h0000;
      coeffs_in_data_log_force[4116] <= 16'h0000;
      coeffs_in_data_log_force[4117] <= 16'h0000;
      coeffs_in_data_log_force[4118] <= 16'h0000;
      coeffs_in_data_log_force[4119] <= 16'h0000;
      coeffs_in_data_log_force[4120] <= 16'h0000;
      coeffs_in_data_log_force[4121] <= 16'h0000;
      coeffs_in_data_log_force[4122] <= 16'h0000;
      coeffs_in_data_log_force[4123] <= 16'h0000;
      coeffs_in_data_log_force[4124] <= 16'h0000;
      coeffs_in_data_log_force[4125] <= 16'h0000;
      coeffs_in_data_log_force[4126] <= 16'h0000;
      coeffs_in_data_log_force[4127] <= 16'h0000;
      coeffs_in_data_log_force[4128] <= 16'h0000;
      coeffs_in_data_log_force[4129] <= 16'h0000;
      coeffs_in_data_log_force[4130] <= 16'h0000;
      coeffs_in_data_log_force[4131] <= 16'h0000;
      coeffs_in_data_log_force[4132] <= 16'h0000;
      coeffs_in_data_log_force[4133] <= 16'h0000;
      coeffs_in_data_log_force[4134] <= 16'h0000;
      coeffs_in_data_log_force[4135] <= 16'h0000;
      coeffs_in_data_log_force[4136] <= 16'h0000;
      coeffs_in_data_log_force[4137] <= 16'h0000;
      coeffs_in_data_log_force[4138] <= 16'h0000;
      coeffs_in_data_log_force[4139] <= 16'h0000;
      coeffs_in_data_log_force[4140] <= 16'h0000;
      coeffs_in_data_log_force[4141] <= 16'h0000;
      coeffs_in_data_log_force[4142] <= 16'h0000;
      coeffs_in_data_log_force[4143] <= 16'h0000;
      coeffs_in_data_log_force[4144] <= 16'h0000;
      coeffs_in_data_log_force[4145] <= 16'h0000;
      coeffs_in_data_log_force[4146] <= 16'h0000;
      coeffs_in_data_log_force[4147] <= 16'h0000;
      coeffs_in_data_log_force[4148] <= 16'h0000;
      coeffs_in_data_log_force[4149] <= 16'h0000;
      coeffs_in_data_log_force[4150] <= 16'h0000;
      coeffs_in_data_log_force[4151] <= 16'h0000;
      coeffs_in_data_log_force[4152] <= 16'h0000;
      coeffs_in_data_log_force[4153] <= 16'h0000;
      coeffs_in_data_log_force[4154] <= 16'h0000;
      coeffs_in_data_log_force[4155] <= 16'h0000;
      coeffs_in_data_log_force[4156] <= 16'h0000;
      coeffs_in_data_log_force[4157] <= 16'h0000;
      coeffs_in_data_log_force[4158] <= 16'h0000;
      coeffs_in_data_log_force[4159] <= 16'h0000;
      coeffs_in_data_log_force[4160] <= 16'h0000;
      coeffs_in_data_log_force[4161] <= 16'h0000;
      coeffs_in_data_log_force[4162] <= 16'h0000;
      coeffs_in_data_log_force[4163] <= 16'h0000;
      coeffs_in_data_log_force[4164] <= 16'h0000;
      coeffs_in_data_log_force[4165] <= 16'h0000;
      coeffs_in_data_log_force[4166] <= 16'h0000;
      coeffs_in_data_log_force[4167] <= 16'h0000;
      coeffs_in_data_log_force[4168] <= 16'h0000;
      coeffs_in_data_log_force[4169] <= 16'h0000;
      coeffs_in_data_log_force[4170] <= 16'h0000;
      coeffs_in_data_log_force[4171] <= 16'h0000;
      coeffs_in_data_log_force[4172] <= 16'h0000;
      coeffs_in_data_log_force[4173] <= 16'h0000;
      coeffs_in_data_log_force[4174] <= 16'h0000;
      coeffs_in_data_log_force[4175] <= 16'h0000;
      coeffs_in_data_log_force[4176] <= 16'h0000;
      coeffs_in_data_log_force[4177] <= 16'h0000;
      coeffs_in_data_log_force[4178] <= 16'h0000;
      coeffs_in_data_log_force[4179] <= 16'h0000;
      coeffs_in_data_log_force[4180] <= 16'h0000;
      coeffs_in_data_log_force[4181] <= 16'h0000;
      coeffs_in_data_log_force[4182] <= 16'h0000;
      coeffs_in_data_log_force[4183] <= 16'h0000;
      coeffs_in_data_log_force[4184] <= 16'h0000;
      coeffs_in_data_log_force[4185] <= 16'h0000;
      coeffs_in_data_log_force[4186] <= 16'h0000;
      coeffs_in_data_log_force[4187] <= 16'h0000;
      coeffs_in_data_log_force[4188] <= 16'h0000;
      coeffs_in_data_log_force[4189] <= 16'h0000;
      coeffs_in_data_log_force[4190] <= 16'h0000;
      coeffs_in_data_log_force[4191] <= 16'h0000;
      coeffs_in_data_log_force[4192] <= 16'h0000;
      coeffs_in_data_log_force[4193] <= 16'h0000;
      coeffs_in_data_log_force[4194] <= 16'h0000;
      coeffs_in_data_log_force[4195] <= 16'h0000;
      coeffs_in_data_log_force[4196] <= 16'h0000;
      coeffs_in_data_log_force[4197] <= 16'h0000;
      coeffs_in_data_log_force[4198] <= 16'h0000;
      coeffs_in_data_log_force[4199] <= 16'h0000;
      coeffs_in_data_log_force[4200] <= 16'h0000;
      coeffs_in_data_log_force[4201] <= 16'h0000;
      coeffs_in_data_log_force[4202] <= 16'h0000;
      coeffs_in_data_log_force[4203] <= 16'h0000;
      coeffs_in_data_log_force[4204] <= 16'h0000;
      coeffs_in_data_log_force[4205] <= 16'h0000;
      coeffs_in_data_log_force[4206] <= 16'h0000;
      coeffs_in_data_log_force[4207] <= 16'h0000;
      coeffs_in_data_log_force[4208] <= 16'h0000;
      coeffs_in_data_log_force[4209] <= 16'h0000;
      coeffs_in_data_log_force[4210] <= 16'h0000;
      coeffs_in_data_log_force[4211] <= 16'h0000;
      coeffs_in_data_log_force[4212] <= 16'h0000;
      coeffs_in_data_log_force[4213] <= 16'h0000;
      coeffs_in_data_log_force[4214] <= 16'h0000;
      coeffs_in_data_log_force[4215] <= 16'h0000;
      coeffs_in_data_log_force[4216] <= 16'h0000;
      coeffs_in_data_log_force[4217] <= 16'h0000;
      coeffs_in_data_log_force[4218] <= 16'h0000;
      coeffs_in_data_log_force[4219] <= 16'h0000;
      coeffs_in_data_log_force[4220] <= 16'h0000;
      coeffs_in_data_log_force[4221] <= 16'h0000;
      coeffs_in_data_log_force[4222] <= 16'h0000;
      coeffs_in_data_log_force[4223] <= 16'h0000;
      coeffs_in_data_log_force[4224] <= 16'h0000;
      coeffs_in_data_log_force[4225] <= 16'h0000;
      coeffs_in_data_log_force[4226] <= 16'h0000;
      coeffs_in_data_log_force[4227] <= 16'h0000;
      coeffs_in_data_log_force[4228] <= 16'h0000;
      coeffs_in_data_log_force[4229] <= 16'h0000;
      coeffs_in_data_log_force[4230] <= 16'h0000;
      coeffs_in_data_log_force[4231] <= 16'h0000;
      coeffs_in_data_log_force[4232] <= 16'h0000;
      coeffs_in_data_log_force[4233] <= 16'h0000;
      coeffs_in_data_log_force[4234] <= 16'h0000;
      coeffs_in_data_log_force[4235] <= 16'h0000;
      coeffs_in_data_log_force[4236] <= 16'h0000;
      coeffs_in_data_log_force[4237] <= 16'h0000;
      coeffs_in_data_log_force[4238] <= 16'h0000;
      coeffs_in_data_log_force[4239] <= 16'h0000;
      coeffs_in_data_log_force[4240] <= 16'h0000;
      coeffs_in_data_log_force[4241] <= 16'h0000;
      coeffs_in_data_log_force[4242] <= 16'h0000;
      coeffs_in_data_log_force[4243] <= 16'h0000;
      coeffs_in_data_log_force[4244] <= 16'h0000;
      coeffs_in_data_log_force[4245] <= 16'h0000;
      coeffs_in_data_log_force[4246] <= 16'h0000;
      coeffs_in_data_log_force[4247] <= 16'h0000;
      coeffs_in_data_log_force[4248] <= 16'h0000;
      coeffs_in_data_log_force[4249] <= 16'h0000;
      coeffs_in_data_log_force[4250] <= 16'h0000;
      coeffs_in_data_log_force[4251] <= 16'h0000;
      coeffs_in_data_log_force[4252] <= 16'h0000;
      coeffs_in_data_log_force[4253] <= 16'h0000;
      coeffs_in_data_log_force[4254] <= 16'h0000;
      coeffs_in_data_log_force[4255] <= 16'h0000;
      coeffs_in_data_log_force[4256] <= 16'h0000;
      coeffs_in_data_log_force[4257] <= 16'h0000;
      coeffs_in_data_log_force[4258] <= 16'h0000;
      coeffs_in_data_log_force[4259] <= 16'h0000;
      coeffs_in_data_log_force[4260] <= 16'h0000;
      coeffs_in_data_log_force[4261] <= 16'h0000;
      coeffs_in_data_log_force[4262] <= 16'h0000;
      coeffs_in_data_log_force[4263] <= 16'h0000;
      coeffs_in_data_log_force[4264] <= 16'h0000;
      coeffs_in_data_log_force[4265] <= 16'h0000;
      coeffs_in_data_log_force[4266] <= 16'h0000;
      coeffs_in_data_log_force[4267] <= 16'h0000;
      coeffs_in_data_log_force[4268] <= 16'h0000;
      coeffs_in_data_log_force[4269] <= 16'h0000;
      coeffs_in_data_log_force[4270] <= 16'h0000;
      coeffs_in_data_log_force[4271] <= 16'h0000;
      coeffs_in_data_log_force[4272] <= 16'h0000;
      coeffs_in_data_log_force[4273] <= 16'h0000;
      coeffs_in_data_log_force[4274] <= 16'h0000;
      coeffs_in_data_log_force[4275] <= 16'h0000;
      coeffs_in_data_log_force[4276] <= 16'h0000;
      coeffs_in_data_log_force[4277] <= 16'h0000;
      coeffs_in_data_log_force[4278] <= 16'h0000;
      coeffs_in_data_log_force[4279] <= 16'h0000;
      coeffs_in_data_log_force[4280] <= 16'h0000;
      coeffs_in_data_log_force[4281] <= 16'h0000;
      coeffs_in_data_log_force[4282] <= 16'h0000;
      coeffs_in_data_log_force[4283] <= 16'h0000;
      coeffs_in_data_log_force[4284] <= 16'h0000;
      coeffs_in_data_log_force[4285] <= 16'h0000;
      coeffs_in_data_log_force[4286] <= 16'h0000;
      coeffs_in_data_log_force[4287] <= 16'h0000;
      coeffs_in_data_log_force[4288] <= 16'h0000;
      coeffs_in_data_log_force[4289] <= 16'h0000;
      coeffs_in_data_log_force[4290] <= 16'h0000;
      coeffs_in_data_log_force[4291] <= 16'h0000;
      coeffs_in_data_log_force[4292] <= 16'h0000;
      coeffs_in_data_log_force[4293] <= 16'h0000;
      coeffs_in_data_log_force[4294] <= 16'h0000;
      coeffs_in_data_log_force[4295] <= 16'h0000;
      coeffs_in_data_log_force[4296] <= 16'h0000;
      coeffs_in_data_log_force[4297] <= 16'h0000;
      coeffs_in_data_log_force[4298] <= 16'h0000;
      coeffs_in_data_log_force[4299] <= 16'h0000;
      coeffs_in_data_log_force[4300] <= 16'h0000;
      coeffs_in_data_log_force[4301] <= 16'h0000;
      coeffs_in_data_log_force[4302] <= 16'h0000;
      coeffs_in_data_log_force[4303] <= 16'h0000;
      coeffs_in_data_log_force[4304] <= 16'h0000;
      coeffs_in_data_log_force[4305] <= 16'h0000;
      coeffs_in_data_log_force[4306] <= 16'h0000;
      coeffs_in_data_log_force[4307] <= 16'h0000;
      coeffs_in_data_log_force[4308] <= 16'h0000;
      coeffs_in_data_log_force[4309] <= 16'h0000;
      coeffs_in_data_log_force[4310] <= 16'h0000;
      coeffs_in_data_log_force[4311] <= 16'h0000;
      coeffs_in_data_log_force[4312] <= 16'h0000;
      coeffs_in_data_log_force[4313] <= 16'h0000;
      coeffs_in_data_log_force[4314] <= 16'h0000;
      coeffs_in_data_log_force[4315] <= 16'h0000;
      coeffs_in_data_log_force[4316] <= 16'h0000;
      coeffs_in_data_log_force[4317] <= 16'h0000;
      coeffs_in_data_log_force[4318] <= 16'h0000;
      coeffs_in_data_log_force[4319] <= 16'h0000;
      coeffs_in_data_log_force[4320] <= 16'h0000;
      coeffs_in_data_log_force[4321] <= 16'h0000;
      coeffs_in_data_log_force[4322] <= 16'h0000;
      coeffs_in_data_log_force[4323] <= 16'h0000;
      coeffs_in_data_log_force[4324] <= 16'h0000;
      coeffs_in_data_log_force[4325] <= 16'h0000;
      coeffs_in_data_log_force[4326] <= 16'h0000;
      coeffs_in_data_log_force[4327] <= 16'h0000;
      coeffs_in_data_log_force[4328] <= 16'h0000;
      coeffs_in_data_log_force[4329] <= 16'h0000;
      coeffs_in_data_log_force[4330] <= 16'h0000;
      coeffs_in_data_log_force[4331] <= 16'h0000;
      coeffs_in_data_log_force[4332] <= 16'h0000;
      coeffs_in_data_log_force[4333] <= 16'h0000;
      coeffs_in_data_log_force[4334] <= 16'h0000;
      coeffs_in_data_log_force[4335] <= 16'h0000;
      coeffs_in_data_log_force[4336] <= 16'h0000;
      coeffs_in_data_log_force[4337] <= 16'h0000;
      coeffs_in_data_log_force[4338] <= 16'h0000;
      coeffs_in_data_log_force[4339] <= 16'h0000;
      coeffs_in_data_log_force[4340] <= 16'h0000;
      coeffs_in_data_log_force[4341] <= 16'h0000;
      coeffs_in_data_log_force[4342] <= 16'h0000;
      coeffs_in_data_log_force[4343] <= 16'h0000;
      coeffs_in_data_log_force[4344] <= 16'h0000;
      coeffs_in_data_log_force[4345] <= 16'h0000;
      coeffs_in_data_log_force[4346] <= 16'h0000;
      coeffs_in_data_log_force[4347] <= 16'h0000;
      coeffs_in_data_log_force[4348] <= 16'h0000;
      coeffs_in_data_log_force[4349] <= 16'h0000;
      coeffs_in_data_log_force[4350] <= 16'h0000;
      coeffs_in_data_log_force[4351] <= 16'h0000;
      coeffs_in_data_log_force[4352] <= 16'h0000;
      coeffs_in_data_log_force[4353] <= 16'h0000;
      coeffs_in_data_log_force[4354] <= 16'h0000;
      coeffs_in_data_log_force[4355] <= 16'h0000;
      coeffs_in_data_log_force[4356] <= 16'h0000;
      coeffs_in_data_log_force[4357] <= 16'h0000;
      coeffs_in_data_log_force[4358] <= 16'h0000;
      coeffs_in_data_log_force[4359] <= 16'h0000;
      coeffs_in_data_log_force[4360] <= 16'h0000;
      coeffs_in_data_log_force[4361] <= 16'h0000;
      coeffs_in_data_log_force[4362] <= 16'h0000;
      coeffs_in_data_log_force[4363] <= 16'h0000;
      coeffs_in_data_log_force[4364] <= 16'h0000;
      coeffs_in_data_log_force[4365] <= 16'h0000;
      coeffs_in_data_log_force[4366] <= 16'h0000;
      coeffs_in_data_log_force[4367] <= 16'h0000;
      coeffs_in_data_log_force[4368] <= 16'h0000;
      coeffs_in_data_log_force[4369] <= 16'h0000;
      coeffs_in_data_log_force[4370] <= 16'h0000;
      coeffs_in_data_log_force[4371] <= 16'h0000;
      coeffs_in_data_log_force[4372] <= 16'h0000;
      coeffs_in_data_log_force[4373] <= 16'h0000;
      coeffs_in_data_log_force[4374] <= 16'h0000;
      coeffs_in_data_log_force[4375] <= 16'h0000;
      coeffs_in_data_log_force[4376] <= 16'h0000;
      coeffs_in_data_log_force[4377] <= 16'h0000;
      coeffs_in_data_log_force[4378] <= 16'h0000;
      coeffs_in_data_log_force[4379] <= 16'h0000;
      coeffs_in_data_log_force[4380] <= 16'h0000;
      coeffs_in_data_log_force[4381] <= 16'h0000;
      coeffs_in_data_log_force[4382] <= 16'h0000;
      coeffs_in_data_log_force[4383] <= 16'h0000;
      coeffs_in_data_log_force[4384] <= 16'h0000;
      coeffs_in_data_log_force[4385] <= 16'h0000;
      coeffs_in_data_log_force[4386] <= 16'h0000;
      coeffs_in_data_log_force[4387] <= 16'h0000;
      coeffs_in_data_log_force[4388] <= 16'h0000;
      coeffs_in_data_log_force[4389] <= 16'h0000;
      coeffs_in_data_log_force[4390] <= 16'h0000;
      coeffs_in_data_log_force[4391] <= 16'h0000;
      coeffs_in_data_log_force[4392] <= 16'h0000;
      coeffs_in_data_log_force[4393] <= 16'h0000;
      coeffs_in_data_log_force[4394] <= 16'h0000;
      coeffs_in_data_log_force[4395] <= 16'h0000;
      coeffs_in_data_log_force[4396] <= 16'h0000;
      coeffs_in_data_log_force[4397] <= 16'h0000;
      coeffs_in_data_log_force[4398] <= 16'h0000;
      coeffs_in_data_log_force[4399] <= 16'h0000;
      coeffs_in_data_log_force[4400] <= 16'h0000;
      coeffs_in_data_log_force[4401] <= 16'h0000;
      coeffs_in_data_log_force[4402] <= 16'h0000;
      coeffs_in_data_log_force[4403] <= 16'h0000;
      coeffs_in_data_log_force[4404] <= 16'h0000;
      coeffs_in_data_log_force[4405] <= 16'h0000;
      coeffs_in_data_log_force[4406] <= 16'h0000;
      coeffs_in_data_log_force[4407] <= 16'h0000;
      coeffs_in_data_log_force[4408] <= 16'h0000;
      coeffs_in_data_log_force[4409] <= 16'h0000;
      coeffs_in_data_log_force[4410] <= 16'h0000;
      coeffs_in_data_log_force[4411] <= 16'h0000;
      coeffs_in_data_log_force[4412] <= 16'h0000;
      coeffs_in_data_log_force[4413] <= 16'h0000;
      coeffs_in_data_log_force[4414] <= 16'h0000;
      coeffs_in_data_log_force[4415] <= 16'h0000;
      coeffs_in_data_log_force[4416] <= 16'h0000;
      coeffs_in_data_log_force[4417] <= 16'h0000;
      coeffs_in_data_log_force[4418] <= 16'h0000;
      coeffs_in_data_log_force[4419] <= 16'h0000;
      coeffs_in_data_log_force[4420] <= 16'h0000;
      coeffs_in_data_log_force[4421] <= 16'h0000;
      coeffs_in_data_log_force[4422] <= 16'h0000;
      coeffs_in_data_log_force[4423] <= 16'h0000;
      coeffs_in_data_log_force[4424] <= 16'h0000;
      coeffs_in_data_log_force[4425] <= 16'h0000;
      coeffs_in_data_log_force[4426] <= 16'h0000;
      coeffs_in_data_log_force[4427] <= 16'h0000;
      coeffs_in_data_log_force[4428] <= 16'h0000;
      coeffs_in_data_log_force[4429] <= 16'h0000;
      coeffs_in_data_log_force[4430] <= 16'h0000;
      coeffs_in_data_log_force[4431] <= 16'h0000;
      coeffs_in_data_log_force[4432] <= 16'h0000;
      coeffs_in_data_log_force[4433] <= 16'h0000;
      coeffs_in_data_log_force[4434] <= 16'h0000;
      coeffs_in_data_log_force[4435] <= 16'h0000;
      coeffs_in_data_log_force[4436] <= 16'h0000;
      coeffs_in_data_log_force[4437] <= 16'h0000;
      coeffs_in_data_log_force[4438] <= 16'h0000;
      coeffs_in_data_log_force[4439] <= 16'h0000;
      coeffs_in_data_log_force[4440] <= 16'h0000;
      coeffs_in_data_log_force[4441] <= 16'h0000;
      coeffs_in_data_log_force[4442] <= 16'h0000;
      coeffs_in_data_log_force[4443] <= 16'h0000;
      coeffs_in_data_log_force[4444] <= 16'h0000;
      coeffs_in_data_log_force[4445] <= 16'h0000;
      coeffs_in_data_log_force[4446] <= 16'h0000;
      coeffs_in_data_log_force[4447] <= 16'h0000;
      coeffs_in_data_log_force[4448] <= 16'h0000;
      coeffs_in_data_log_force[4449] <= 16'h0000;
      coeffs_in_data_log_force[4450] <= 16'h0000;
      coeffs_in_data_log_force[4451] <= 16'h0000;
      coeffs_in_data_log_force[4452] <= 16'h0000;
      coeffs_in_data_log_force[4453] <= 16'h0000;
      coeffs_in_data_log_force[4454] <= 16'h0000;
      coeffs_in_data_log_force[4455] <= 16'h0000;
      coeffs_in_data_log_force[4456] <= 16'h0000;
      coeffs_in_data_log_force[4457] <= 16'h0000;
      coeffs_in_data_log_force[4458] <= 16'h0000;
      coeffs_in_data_log_force[4459] <= 16'h0000;
      coeffs_in_data_log_force[4460] <= 16'h0000;
      coeffs_in_data_log_force[4461] <= 16'h0000;
      coeffs_in_data_log_force[4462] <= 16'h0000;
      coeffs_in_data_log_force[4463] <= 16'h0000;
      coeffs_in_data_log_force[4464] <= 16'h0000;
      coeffs_in_data_log_force[4465] <= 16'h0000;
      coeffs_in_data_log_force[4466] <= 16'h0000;
      coeffs_in_data_log_force[4467] <= 16'h0000;
      coeffs_in_data_log_force[4468] <= 16'h0000;
      coeffs_in_data_log_force[4469] <= 16'h0000;
      coeffs_in_data_log_force[4470] <= 16'h0000;
      coeffs_in_data_log_force[4471] <= 16'h0000;
      coeffs_in_data_log_force[4472] <= 16'h0000;
      coeffs_in_data_log_force[4473] <= 16'h0000;
      coeffs_in_data_log_force[4474] <= 16'h0000;
      coeffs_in_data_log_force[4475] <= 16'h0000;
      coeffs_in_data_log_force[4476] <= 16'h0000;
      coeffs_in_data_log_force[4477] <= 16'h0000;
      coeffs_in_data_log_force[4478] <= 16'h0000;
      coeffs_in_data_log_force[4479] <= 16'h0000;
      coeffs_in_data_log_force[4480] <= 16'h0000;
      coeffs_in_data_log_force[4481] <= 16'h0000;
      coeffs_in_data_log_force[4482] <= 16'h0000;
      coeffs_in_data_log_force[4483] <= 16'h0000;
      coeffs_in_data_log_force[4484] <= 16'h0000;
      coeffs_in_data_log_force[4485] <= 16'h0000;
      coeffs_in_data_log_force[4486] <= 16'h0000;
      coeffs_in_data_log_force[4487] <= 16'h0000;
      coeffs_in_data_log_force[4488] <= 16'h0000;
      coeffs_in_data_log_force[4489] <= 16'h0000;
      coeffs_in_data_log_force[4490] <= 16'h0000;
      coeffs_in_data_log_force[4491] <= 16'h0000;
      coeffs_in_data_log_force[4492] <= 16'h0000;
      coeffs_in_data_log_force[4493] <= 16'h0000;
      coeffs_in_data_log_force[4494] <= 16'h0000;
      coeffs_in_data_log_force[4495] <= 16'h0000;
      coeffs_in_data_log_force[4496] <= 16'h0000;
      coeffs_in_data_log_force[4497] <= 16'h0000;
      coeffs_in_data_log_force[4498] <= 16'h0000;
      coeffs_in_data_log_force[4499] <= 16'h0000;
      coeffs_in_data_log_force[4500] <= 16'h0000;
      coeffs_in_data_log_force[4501] <= 16'h0000;
      coeffs_in_data_log_force[4502] <= 16'h0000;
      coeffs_in_data_log_force[4503] <= 16'h0000;
      coeffs_in_data_log_force[4504] <= 16'h0000;
      coeffs_in_data_log_force[4505] <= 16'h0000;
      coeffs_in_data_log_force[4506] <= 16'h0000;
      coeffs_in_data_log_force[4507] <= 16'h0000;
      coeffs_in_data_log_force[4508] <= 16'h0000;
      coeffs_in_data_log_force[4509] <= 16'h0000;
      coeffs_in_data_log_force[4510] <= 16'h0000;
      coeffs_in_data_log_force[4511] <= 16'h0000;
      coeffs_in_data_log_force[4512] <= 16'h0000;
      coeffs_in_data_log_force[4513] <= 16'h0000;
      coeffs_in_data_log_force[4514] <= 16'h0000;
      coeffs_in_data_log_force[4515] <= 16'h0000;
      coeffs_in_data_log_force[4516] <= 16'h0000;
      coeffs_in_data_log_force[4517] <= 16'h0000;
      coeffs_in_data_log_force[4518] <= 16'h0000;
      coeffs_in_data_log_force[4519] <= 16'h0000;
      coeffs_in_data_log_force[4520] <= 16'h0000;
      coeffs_in_data_log_force[4521] <= 16'h0000;
      coeffs_in_data_log_force[4522] <= 16'h0000;
      coeffs_in_data_log_force[4523] <= 16'h0000;
      coeffs_in_data_log_force[4524] <= 16'h0000;
      coeffs_in_data_log_force[4525] <= 16'h0000;
      coeffs_in_data_log_force[4526] <= 16'h0000;
      coeffs_in_data_log_force[4527] <= 16'h0000;
      coeffs_in_data_log_force[4528] <= 16'h0000;
      coeffs_in_data_log_force[4529] <= 16'h0000;
      coeffs_in_data_log_force[4530] <= 16'h0000;
      coeffs_in_data_log_force[4531] <= 16'h0000;
      coeffs_in_data_log_force[4532] <= 16'h0000;
      coeffs_in_data_log_force[4533] <= 16'h0000;
      coeffs_in_data_log_force[4534] <= 16'h0000;
      coeffs_in_data_log_force[4535] <= 16'h0000;
      coeffs_in_data_log_force[4536] <= 16'h0000;
      coeffs_in_data_log_force[4537] <= 16'h0000;
      coeffs_in_data_log_force[4538] <= 16'h0000;
      coeffs_in_data_log_force[4539] <= 16'h0000;
      coeffs_in_data_log_force[4540] <= 16'h0000;
      coeffs_in_data_log_force[4541] <= 16'h0000;
      coeffs_in_data_log_force[4542] <= 16'h0000;
      coeffs_in_data_log_force[4543] <= 16'h0000;
      coeffs_in_data_log_force[4544] <= 16'h0000;
      coeffs_in_data_log_force[4545] <= 16'h0000;
      coeffs_in_data_log_force[4546] <= 16'h0000;
      coeffs_in_data_log_force[4547] <= 16'h0000;
      coeffs_in_data_log_force[4548] <= 16'h0000;
      coeffs_in_data_log_force[4549] <= 16'h0000;
      coeffs_in_data_log_force[4550] <= 16'h0000;
      coeffs_in_data_log_force[4551] <= 16'h0000;
      coeffs_in_data_log_force[4552] <= 16'h0000;
      coeffs_in_data_log_force[4553] <= 16'h0000;
      coeffs_in_data_log_force[4554] <= 16'h0000;
      coeffs_in_data_log_force[4555] <= 16'h0000;
      coeffs_in_data_log_force[4556] <= 16'h0000;
      coeffs_in_data_log_force[4557] <= 16'h0000;
      coeffs_in_data_log_force[4558] <= 16'h0000;
      coeffs_in_data_log_force[4559] <= 16'h0000;
      coeffs_in_data_log_force[4560] <= 16'h0000;
      coeffs_in_data_log_force[4561] <= 16'h0000;
      coeffs_in_data_log_force[4562] <= 16'h0000;
      coeffs_in_data_log_force[4563] <= 16'h0000;
      coeffs_in_data_log_force[4564] <= 16'h0000;
      coeffs_in_data_log_force[4565] <= 16'h0000;
      coeffs_in_data_log_force[4566] <= 16'h0000;
      coeffs_in_data_log_force[4567] <= 16'h0000;
      coeffs_in_data_log_force[4568] <= 16'h0000;
      coeffs_in_data_log_force[4569] <= 16'h0000;
      coeffs_in_data_log_force[4570] <= 16'h0000;
      coeffs_in_data_log_force[4571] <= 16'h0000;
      coeffs_in_data_log_force[4572] <= 16'h0000;
      coeffs_in_data_log_force[4573] <= 16'h0000;
      coeffs_in_data_log_force[4574] <= 16'h0000;
      coeffs_in_data_log_force[4575] <= 16'h0000;
      coeffs_in_data_log_force[4576] <= 16'h0000;
      coeffs_in_data_log_force[4577] <= 16'h0000;
      coeffs_in_data_log_force[4578] <= 16'h0000;
      coeffs_in_data_log_force[4579] <= 16'h0000;
      coeffs_in_data_log_force[4580] <= 16'h0000;
      coeffs_in_data_log_force[4581] <= 16'h0000;
      coeffs_in_data_log_force[4582] <= 16'h0000;
      coeffs_in_data_log_force[4583] <= 16'h0000;
      coeffs_in_data_log_force[4584] <= 16'h0000;
      coeffs_in_data_log_force[4585] <= 16'h0000;
      coeffs_in_data_log_force[4586] <= 16'h0000;
      coeffs_in_data_log_force[4587] <= 16'h0000;
      coeffs_in_data_log_force[4588] <= 16'h0000;
      coeffs_in_data_log_force[4589] <= 16'h0000;
      coeffs_in_data_log_force[4590] <= 16'h0000;
      coeffs_in_data_log_force[4591] <= 16'h0000;
      coeffs_in_data_log_force[4592] <= 16'h0000;
      coeffs_in_data_log_force[4593] <= 16'h0000;
      coeffs_in_data_log_force[4594] <= 16'h0000;
      coeffs_in_data_log_force[4595] <= 16'h0000;
      coeffs_in_data_log_force[4596] <= 16'h0000;
      coeffs_in_data_log_force[4597] <= 16'h0000;
      coeffs_in_data_log_force[4598] <= 16'h0000;
      coeffs_in_data_log_force[4599] <= 16'h0000;
      coeffs_in_data_log_force[4600] <= 16'h0000;
      coeffs_in_data_log_force[4601] <= 16'h0000;
      coeffs_in_data_log_force[4602] <= 16'h0000;
      coeffs_in_data_log_force[4603] <= 16'h0000;
      coeffs_in_data_log_force[4604] <= 16'h0000;
      coeffs_in_data_log_force[4605] <= 16'h0000;
      coeffs_in_data_log_force[4606] <= 16'h0000;
      coeffs_in_data_log_force[4607] <= 16'h0000;
      coeffs_in_data_log_force[4608] <= 16'h0000;
      coeffs_in_data_log_force[4609] <= 16'h0000;
      coeffs_in_data_log_force[4610] <= 16'h0000;
      coeffs_in_data_log_force[4611] <= 16'h0000;
      coeffs_in_data_log_force[4612] <= 16'h0000;
      coeffs_in_data_log_force[4613] <= 16'h0000;
      coeffs_in_data_log_force[4614] <= 16'h0000;
      coeffs_in_data_log_force[4615] <= 16'h0000;
      coeffs_in_data_log_force[4616] <= 16'h0000;
      coeffs_in_data_log_force[4617] <= 16'h0000;
      coeffs_in_data_log_force[4618] <= 16'h0000;
      coeffs_in_data_log_force[4619] <= 16'h0000;
      coeffs_in_data_log_force[4620] <= 16'h0000;
      coeffs_in_data_log_force[4621] <= 16'h0000;
      coeffs_in_data_log_force[4622] <= 16'h0000;
      coeffs_in_data_log_force[4623] <= 16'h0000;
      coeffs_in_data_log_force[4624] <= 16'h0000;
      coeffs_in_data_log_force[4625] <= 16'h0000;
      coeffs_in_data_log_force[4626] <= 16'h0000;
      coeffs_in_data_log_force[4627] <= 16'h0000;
      coeffs_in_data_log_force[4628] <= 16'h0000;
      coeffs_in_data_log_force[4629] <= 16'h0000;
      coeffs_in_data_log_force[4630] <= 16'h0000;
      coeffs_in_data_log_force[4631] <= 16'h0000;
      coeffs_in_data_log_force[4632] <= 16'h0000;
      coeffs_in_data_log_force[4633] <= 16'h0000;
      coeffs_in_data_log_force[4634] <= 16'h0000;
      coeffs_in_data_log_force[4635] <= 16'h0000;
      coeffs_in_data_log_force[4636] <= 16'h0000;
      coeffs_in_data_log_force[4637] <= 16'h0000;
      coeffs_in_data_log_force[4638] <= 16'h0000;
      coeffs_in_data_log_force[4639] <= 16'h0000;
      coeffs_in_data_log_force[4640] <= 16'h0000;
      coeffs_in_data_log_force[4641] <= 16'h0000;
      coeffs_in_data_log_force[4642] <= 16'h0000;
      coeffs_in_data_log_force[4643] <= 16'h0000;
      coeffs_in_data_log_force[4644] <= 16'h0000;
      coeffs_in_data_log_force[4645] <= 16'h0000;
      coeffs_in_data_log_force[4646] <= 16'h0000;
      coeffs_in_data_log_force[4647] <= 16'h0000;
      coeffs_in_data_log_force[4648] <= 16'h0000;
      coeffs_in_data_log_force[4649] <= 16'h0000;
      coeffs_in_data_log_force[4650] <= 16'h0000;
      coeffs_in_data_log_force[4651] <= 16'h0000;
      coeffs_in_data_log_force[4652] <= 16'h0000;
      coeffs_in_data_log_force[4653] <= 16'h0000;
      coeffs_in_data_log_force[4654] <= 16'h0000;
      coeffs_in_data_log_force[4655] <= 16'h0000;
      coeffs_in_data_log_force[4656] <= 16'h0000;
      coeffs_in_data_log_force[4657] <= 16'h0000;
      coeffs_in_data_log_force[4658] <= 16'h0000;
      coeffs_in_data_log_force[4659] <= 16'h0000;
      coeffs_in_data_log_force[4660] <= 16'h0000;
      coeffs_in_data_log_force[4661] <= 16'h0000;
      coeffs_in_data_log_force[4662] <= 16'h0000;
      coeffs_in_data_log_force[4663] <= 16'h0000;
      coeffs_in_data_log_force[4664] <= 16'h0000;
      coeffs_in_data_log_force[4665] <= 16'h0000;
      coeffs_in_data_log_force[4666] <= 16'h0000;
      coeffs_in_data_log_force[4667] <= 16'h0000;
      coeffs_in_data_log_force[4668] <= 16'h0000;
      coeffs_in_data_log_force[4669] <= 16'h0000;
      coeffs_in_data_log_force[4670] <= 16'h0000;
      coeffs_in_data_log_force[4671] <= 16'h0000;
      coeffs_in_data_log_force[4672] <= 16'h0000;
      coeffs_in_data_log_force[4673] <= 16'h0000;
      coeffs_in_data_log_force[4674] <= 16'h0000;
      coeffs_in_data_log_force[4675] <= 16'h0000;
      coeffs_in_data_log_force[4676] <= 16'h0000;
      coeffs_in_data_log_force[4677] <= 16'h0000;
      coeffs_in_data_log_force[4678] <= 16'h0000;
      coeffs_in_data_log_force[4679] <= 16'h0000;
      coeffs_in_data_log_force[4680] <= 16'h0000;
      coeffs_in_data_log_force[4681] <= 16'h0000;
      coeffs_in_data_log_force[4682] <= 16'h0000;
      coeffs_in_data_log_force[4683] <= 16'h0000;
      coeffs_in_data_log_force[4684] <= 16'h0000;
      coeffs_in_data_log_force[4685] <= 16'h0000;
      coeffs_in_data_log_force[4686] <= 16'h0000;
      coeffs_in_data_log_force[4687] <= 16'h0000;
      coeffs_in_data_log_force[4688] <= 16'h0000;
      coeffs_in_data_log_force[4689] <= 16'h0000;
      coeffs_in_data_log_force[4690] <= 16'h0000;
      coeffs_in_data_log_force[4691] <= 16'h0000;
      coeffs_in_data_log_force[4692] <= 16'h0000;
      coeffs_in_data_log_force[4693] <= 16'h0000;
      coeffs_in_data_log_force[4694] <= 16'h0000;
      coeffs_in_data_log_force[4695] <= 16'h0000;
      coeffs_in_data_log_force[4696] <= 16'h0000;
      coeffs_in_data_log_force[4697] <= 16'h0000;
      coeffs_in_data_log_force[4698] <= 16'h0000;
      coeffs_in_data_log_force[4699] <= 16'h0000;
      coeffs_in_data_log_force[4700] <= 16'h0000;
      coeffs_in_data_log_force[4701] <= 16'h0000;
      coeffs_in_data_log_force[4702] <= 16'h0000;
      coeffs_in_data_log_force[4703] <= 16'h0000;
      coeffs_in_data_log_force[4704] <= 16'h0000;
      coeffs_in_data_log_force[4705] <= 16'h0000;
      coeffs_in_data_log_force[4706] <= 16'h0000;
      coeffs_in_data_log_force[4707] <= 16'h0000;
      coeffs_in_data_log_force[4708] <= 16'h0000;
      coeffs_in_data_log_force[4709] <= 16'h0000;
      coeffs_in_data_log_force[4710] <= 16'h0000;
      coeffs_in_data_log_force[4711] <= 16'h0000;
      coeffs_in_data_log_force[4712] <= 16'h0000;
      coeffs_in_data_log_force[4713] <= 16'h0000;
      coeffs_in_data_log_force[4714] <= 16'h0000;
      coeffs_in_data_log_force[4715] <= 16'h0000;
      coeffs_in_data_log_force[4716] <= 16'h0000;
      coeffs_in_data_log_force[4717] <= 16'h0000;
      coeffs_in_data_log_force[4718] <= 16'h0000;
      coeffs_in_data_log_force[4719] <= 16'h0000;
      coeffs_in_data_log_force[4720] <= 16'h0000;
      coeffs_in_data_log_force[4721] <= 16'h0000;
      coeffs_in_data_log_force[4722] <= 16'h0000;
      coeffs_in_data_log_force[4723] <= 16'h0000;
      coeffs_in_data_log_force[4724] <= 16'h0000;
      coeffs_in_data_log_force[4725] <= 16'h0000;
      coeffs_in_data_log_force[4726] <= 16'h0000;
      coeffs_in_data_log_force[4727] <= 16'h0000;
      coeffs_in_data_log_force[4728] <= 16'h0000;
      coeffs_in_data_log_force[4729] <= 16'h0000;
      coeffs_in_data_log_force[4730] <= 16'h0000;
      coeffs_in_data_log_force[4731] <= 16'h0000;
      coeffs_in_data_log_force[4732] <= 16'h0000;
      coeffs_in_data_log_force[4733] <= 16'h0000;
      coeffs_in_data_log_force[4734] <= 16'h0000;
      coeffs_in_data_log_force[4735] <= 16'h0000;
      coeffs_in_data_log_force[4736] <= 16'h0000;
      coeffs_in_data_log_force[4737] <= 16'h0000;
      coeffs_in_data_log_force[4738] <= 16'h0000;
      coeffs_in_data_log_force[4739] <= 16'h0000;
      coeffs_in_data_log_force[4740] <= 16'h0000;
      coeffs_in_data_log_force[4741] <= 16'h0000;
      coeffs_in_data_log_force[4742] <= 16'h0000;
      coeffs_in_data_log_force[4743] <= 16'h0000;
      coeffs_in_data_log_force[4744] <= 16'h0000;
      coeffs_in_data_log_force[4745] <= 16'h0000;
      coeffs_in_data_log_force[4746] <= 16'h0000;
      coeffs_in_data_log_force[4747] <= 16'h0000;
      coeffs_in_data_log_force[4748] <= 16'h0000;
      coeffs_in_data_log_force[4749] <= 16'h0000;
      coeffs_in_data_log_force[4750] <= 16'h0000;
      coeffs_in_data_log_force[4751] <= 16'h0000;
      coeffs_in_data_log_force[4752] <= 16'h0000;
      coeffs_in_data_log_force[4753] <= 16'h0000;
      coeffs_in_data_log_force[4754] <= 16'h0000;
      coeffs_in_data_log_force[4755] <= 16'h0000;
      coeffs_in_data_log_force[4756] <= 16'h0000;
      coeffs_in_data_log_force[4757] <= 16'h0000;
      coeffs_in_data_log_force[4758] <= 16'h0000;
      coeffs_in_data_log_force[4759] <= 16'h0000;
      coeffs_in_data_log_force[4760] <= 16'h0000;
      coeffs_in_data_log_force[4761] <= 16'h0000;
      coeffs_in_data_log_force[4762] <= 16'h0000;
      coeffs_in_data_log_force[4763] <= 16'h0000;
      coeffs_in_data_log_force[4764] <= 16'h0000;
      coeffs_in_data_log_force[4765] <= 16'h0000;
      coeffs_in_data_log_force[4766] <= 16'h0000;
      coeffs_in_data_log_force[4767] <= 16'h0000;
      coeffs_in_data_log_force[4768] <= 16'h0000;
      coeffs_in_data_log_force[4769] <= 16'h0000;
      coeffs_in_data_log_force[4770] <= 16'h0000;
      coeffs_in_data_log_force[4771] <= 16'h0000;
      coeffs_in_data_log_force[4772] <= 16'h0000;
      coeffs_in_data_log_force[4773] <= 16'h0000;
      coeffs_in_data_log_force[4774] <= 16'h0000;
      coeffs_in_data_log_force[4775] <= 16'h0000;
      coeffs_in_data_log_force[4776] <= 16'h0000;
      coeffs_in_data_log_force[4777] <= 16'h0000;
      coeffs_in_data_log_force[4778] <= 16'h0000;
      coeffs_in_data_log_force[4779] <= 16'h0000;
      coeffs_in_data_log_force[4780] <= 16'h0000;
      coeffs_in_data_log_force[4781] <= 16'h0000;
      coeffs_in_data_log_force[4782] <= 16'h0000;
      coeffs_in_data_log_force[4783] <= 16'h0000;
      coeffs_in_data_log_force[4784] <= 16'h0000;
      coeffs_in_data_log_force[4785] <= 16'h0000;
      coeffs_in_data_log_force[4786] <= 16'h0000;
      coeffs_in_data_log_force[4787] <= 16'h0000;
      coeffs_in_data_log_force[4788] <= 16'h0000;
      coeffs_in_data_log_force[4789] <= 16'h0000;
      coeffs_in_data_log_force[4790] <= 16'h0000;
      coeffs_in_data_log_force[4791] <= 16'h0000;
      coeffs_in_data_log_force[4792] <= 16'h0000;
      coeffs_in_data_log_force[4793] <= 16'h0000;
      coeffs_in_data_log_force[4794] <= 16'h0000;
      coeffs_in_data_log_force[4795] <= 16'h0000;
      coeffs_in_data_log_force[4796] <= 16'h0000;
      coeffs_in_data_log_force[4797] <= 16'h0000;
      coeffs_in_data_log_force[4798] <= 16'h0000;
      coeffs_in_data_log_force[4799] <= 16'h0000;
      coeffs_in_data_log_force[4800] <= 16'h0000;
      coeffs_in_data_log_force[4801] <= 16'h0000;
      coeffs_in_data_log_force[4802] <= 16'h0000;
      coeffs_in_data_log_force[4803] <= 16'h0000;
      coeffs_in_data_log_force[4804] <= 16'h0000;
      coeffs_in_data_log_force[4805] <= 16'h0000;
      coeffs_in_data_log_force[4806] <= 16'h0000;
      coeffs_in_data_log_force[4807] <= 16'h0000;
      coeffs_in_data_log_force[4808] <= 16'h0000;
      coeffs_in_data_log_force[4809] <= 16'h0000;
      coeffs_in_data_log_force[4810] <= 16'h0000;
      coeffs_in_data_log_force[4811] <= 16'h0000;
      coeffs_in_data_log_force[4812] <= 16'h0000;
      coeffs_in_data_log_force[4813] <= 16'h0000;
      coeffs_in_data_log_force[4814] <= 16'h0000;
      coeffs_in_data_log_force[4815] <= 16'h0000;
      coeffs_in_data_log_force[4816] <= 16'h0000;
      coeffs_in_data_log_force[4817] <= 16'h0000;
      coeffs_in_data_log_force[4818] <= 16'h0000;
      coeffs_in_data_log_force[4819] <= 16'h0000;
      coeffs_in_data_log_force[4820] <= 16'h0000;
      coeffs_in_data_log_force[4821] <= 16'h0000;
      coeffs_in_data_log_force[4822] <= 16'h0000;
      coeffs_in_data_log_force[4823] <= 16'h0000;
      coeffs_in_data_log_force[4824] <= 16'h0000;
      coeffs_in_data_log_force[4825] <= 16'h0000;
      coeffs_in_data_log_force[4826] <= 16'h0000;
      coeffs_in_data_log_force[4827] <= 16'h0000;
      coeffs_in_data_log_force[4828] <= 16'h0000;
      coeffs_in_data_log_force[4829] <= 16'h0000;
      coeffs_in_data_log_force[4830] <= 16'h0000;
      coeffs_in_data_log_force[4831] <= 16'h0000;
      coeffs_in_data_log_force[4832] <= 16'h0000;
      coeffs_in_data_log_force[4833] <= 16'h0000;
      coeffs_in_data_log_force[4834] <= 16'h0000;
      coeffs_in_data_log_force[4835] <= 16'h0000;
      coeffs_in_data_log_force[4836] <= 16'h0000;
      coeffs_in_data_log_force[4837] <= 16'h0000;
      coeffs_in_data_log_force[4838] <= 16'h0000;
      coeffs_in_data_log_force[4839] <= 16'h0000;
      coeffs_in_data_log_force[4840] <= 16'h0000;
      coeffs_in_data_log_force[4841] <= 16'h0000;
      coeffs_in_data_log_force[4842] <= 16'h0000;
      coeffs_in_data_log_force[4843] <= 16'h0000;
      coeffs_in_data_log_force[4844] <= 16'h0000;
      coeffs_in_data_log_force[4845] <= 16'h0000;
      coeffs_in_data_log_force[4846] <= 16'h0000;
      coeffs_in_data_log_force[4847] <= 16'h0000;
      coeffs_in_data_log_force[4848] <= 16'h0000;
      coeffs_in_data_log_force[4849] <= 16'h0000;
      coeffs_in_data_log_force[4850] <= 16'h0000;
      coeffs_in_data_log_force[4851] <= 16'h0000;
      coeffs_in_data_log_force[4852] <= 16'h0000;
      coeffs_in_data_log_force[4853] <= 16'h0000;
      coeffs_in_data_log_force[4854] <= 16'h0000;
      coeffs_in_data_log_force[4855] <= 16'h0000;
      coeffs_in_data_log_force[4856] <= 16'h0000;
      coeffs_in_data_log_force[4857] <= 16'h0000;
      coeffs_in_data_log_force[4858] <= 16'h0000;
      coeffs_in_data_log_force[4859] <= 16'h0000;
      coeffs_in_data_log_force[4860] <= 16'h0000;
      coeffs_in_data_log_force[4861] <= 16'h0000;
      coeffs_in_data_log_force[4862] <= 16'h0000;
      coeffs_in_data_log_force[4863] <= 16'h0000;
      coeffs_in_data_log_force[4864] <= 16'h0000;
      coeffs_in_data_log_force[4865] <= 16'h0000;
      coeffs_in_data_log_force[4866] <= 16'h0000;
      coeffs_in_data_log_force[4867] <= 16'h0000;
      coeffs_in_data_log_force[4868] <= 16'h0000;
      coeffs_in_data_log_force[4869] <= 16'h0000;
      coeffs_in_data_log_force[4870] <= 16'h0000;
      coeffs_in_data_log_force[4871] <= 16'h0000;
      coeffs_in_data_log_force[4872] <= 16'h0000;
      coeffs_in_data_log_force[4873] <= 16'h0000;
      coeffs_in_data_log_force[4874] <= 16'h0000;
      coeffs_in_data_log_force[4875] <= 16'h0000;
      coeffs_in_data_log_force[4876] <= 16'h0000;
      coeffs_in_data_log_force[4877] <= 16'h0000;
      coeffs_in_data_log_force[4878] <= 16'h0000;
      coeffs_in_data_log_force[4879] <= 16'h0000;
      coeffs_in_data_log_force[4880] <= 16'h0000;
      coeffs_in_data_log_force[4881] <= 16'h0000;
      coeffs_in_data_log_force[4882] <= 16'h0000;
      coeffs_in_data_log_force[4883] <= 16'h0000;
      coeffs_in_data_log_force[4884] <= 16'h0000;
      coeffs_in_data_log_force[4885] <= 16'h0000;
      coeffs_in_data_log_force[4886] <= 16'h0000;
      coeffs_in_data_log_force[4887] <= 16'h0000;
      coeffs_in_data_log_force[4888] <= 16'h0000;
      coeffs_in_data_log_force[4889] <= 16'h0000;
      coeffs_in_data_log_force[4890] <= 16'h0000;
      coeffs_in_data_log_force[4891] <= 16'h0000;
      coeffs_in_data_log_force[4892] <= 16'h0000;
      coeffs_in_data_log_force[4893] <= 16'h0000;
      coeffs_in_data_log_force[4894] <= 16'h0000;
      coeffs_in_data_log_force[4895] <= 16'h0000;
      coeffs_in_data_log_force[4896] <= 16'h0000;
      coeffs_in_data_log_force[4897] <= 16'h0000;
      coeffs_in_data_log_force[4898] <= 16'h0000;
      coeffs_in_data_log_force[4899] <= 16'h0000;
      coeffs_in_data_log_force[4900] <= 16'h0000;
      coeffs_in_data_log_force[4901] <= 16'h0000;
      coeffs_in_data_log_force[4902] <= 16'h0000;
      coeffs_in_data_log_force[4903] <= 16'h0000;
      coeffs_in_data_log_force[4904] <= 16'h0000;
      coeffs_in_data_log_force[4905] <= 16'h0000;
      coeffs_in_data_log_force[4906] <= 16'h0000;
      coeffs_in_data_log_force[4907] <= 16'h0000;
      coeffs_in_data_log_force[4908] <= 16'h0000;
      coeffs_in_data_log_force[4909] <= 16'h0000;
      coeffs_in_data_log_force[4910] <= 16'h0000;
      coeffs_in_data_log_force[4911] <= 16'h0000;
      coeffs_in_data_log_force[4912] <= 16'h0000;
      coeffs_in_data_log_force[4913] <= 16'h0000;
      coeffs_in_data_log_force[4914] <= 16'h0000;
      coeffs_in_data_log_force[4915] <= 16'h0000;
      coeffs_in_data_log_force[4916] <= 16'h0000;
      coeffs_in_data_log_force[4917] <= 16'h0000;
      coeffs_in_data_log_force[4918] <= 16'h0000;
      coeffs_in_data_log_force[4919] <= 16'h0000;
      coeffs_in_data_log_force[4920] <= 16'h0000;
      coeffs_in_data_log_force[4921] <= 16'h0000;
      coeffs_in_data_log_force[4922] <= 16'h0000;
      coeffs_in_data_log_force[4923] <= 16'h0000;
      coeffs_in_data_log_force[4924] <= 16'h0000;
      coeffs_in_data_log_force[4925] <= 16'h0000;
      coeffs_in_data_log_force[4926] <= 16'h0000;
      coeffs_in_data_log_force[4927] <= 16'h0000;
      coeffs_in_data_log_force[4928] <= 16'h0000;
      coeffs_in_data_log_force[4929] <= 16'h0000;
      coeffs_in_data_log_force[4930] <= 16'h0000;
      coeffs_in_data_log_force[4931] <= 16'h0000;
      coeffs_in_data_log_force[4932] <= 16'h0000;
      coeffs_in_data_log_force[4933] <= 16'h0000;
      coeffs_in_data_log_force[4934] <= 16'h0000;
      coeffs_in_data_log_force[4935] <= 16'h0000;
      coeffs_in_data_log_force[4936] <= 16'h0000;
      coeffs_in_data_log_force[4937] <= 16'h0000;
      coeffs_in_data_log_force[4938] <= 16'h0000;
      coeffs_in_data_log_force[4939] <= 16'h0000;
      coeffs_in_data_log_force[4940] <= 16'h0000;
      coeffs_in_data_log_force[4941] <= 16'h0000;
      coeffs_in_data_log_force[4942] <= 16'h0000;
      coeffs_in_data_log_force[4943] <= 16'h0000;
      coeffs_in_data_log_force[4944] <= 16'h0000;
      coeffs_in_data_log_force[4945] <= 16'h0000;
      coeffs_in_data_log_force[4946] <= 16'h0000;
      coeffs_in_data_log_force[4947] <= 16'h0000;
      coeffs_in_data_log_force[4948] <= 16'h0000;
      coeffs_in_data_log_force[4949] <= 16'h0000;
      coeffs_in_data_log_force[4950] <= 16'h0000;
      coeffs_in_data_log_force[4951] <= 16'h0000;
      coeffs_in_data_log_force[4952] <= 16'h0000;
      coeffs_in_data_log_force[4953] <= 16'h0000;
      coeffs_in_data_log_force[4954] <= 16'h0000;
      coeffs_in_data_log_force[4955] <= 16'h0000;
      coeffs_in_data_log_force[4956] <= 16'h0000;
      coeffs_in_data_log_force[4957] <= 16'h0000;
      coeffs_in_data_log_force[4958] <= 16'h0000;
      coeffs_in_data_log_force[4959] <= 16'h0000;
      coeffs_in_data_log_force[4960] <= 16'h0000;
      coeffs_in_data_log_force[4961] <= 16'h0000;
      coeffs_in_data_log_force[4962] <= 16'h0000;
      coeffs_in_data_log_force[4963] <= 16'h0000;
      coeffs_in_data_log_force[4964] <= 16'h0000;
      coeffs_in_data_log_force[4965] <= 16'h0000;
      coeffs_in_data_log_force[4966] <= 16'h0000;
      coeffs_in_data_log_force[4967] <= 16'h0000;
      coeffs_in_data_log_force[4968] <= 16'h0000;
      coeffs_in_data_log_force[4969] <= 16'h0000;
      coeffs_in_data_log_force[4970] <= 16'h0000;
      coeffs_in_data_log_force[4971] <= 16'h0000;
      coeffs_in_data_log_force[4972] <= 16'h0000;
      coeffs_in_data_log_force[4973] <= 16'h0000;
      coeffs_in_data_log_force[4974] <= 16'h0000;
      coeffs_in_data_log_force[4975] <= 16'h0000;
      coeffs_in_data_log_force[4976] <= 16'h0000;
      coeffs_in_data_log_force[4977] <= 16'h0000;
      coeffs_in_data_log_force[4978] <= 16'h0000;
      coeffs_in_data_log_force[4979] <= 16'h0000;
      coeffs_in_data_log_force[4980] <= 16'h0000;
      coeffs_in_data_log_force[4981] <= 16'h0000;
      coeffs_in_data_log_force[4982] <= 16'h0000;
      coeffs_in_data_log_force[4983] <= 16'h0000;
      coeffs_in_data_log_force[4984] <= 16'h0000;
      coeffs_in_data_log_force[4985] <= 16'h0000;
      coeffs_in_data_log_force[4986] <= 16'h0000;
      coeffs_in_data_log_force[4987] <= 16'h0000;
      coeffs_in_data_log_force[4988] <= 16'h0000;
      coeffs_in_data_log_force[4989] <= 16'h0000;
      coeffs_in_data_log_force[4990] <= 16'h0000;
      coeffs_in_data_log_force[4991] <= 16'h0000;
      coeffs_in_data_log_force[4992] <= 16'h0000;
      coeffs_in_data_log_force[4993] <= 16'h0000;
      coeffs_in_data_log_force[4994] <= 16'h0000;
      coeffs_in_data_log_force[4995] <= 16'h0000;
      coeffs_in_data_log_force[4996] <= 16'h0000;
      coeffs_in_data_log_force[4997] <= 16'h0000;
      coeffs_in_data_log_force[4998] <= 16'h0000;
      coeffs_in_data_log_force[4999] <= 16'h0000;
      coeffs_in_data_log_force[5000] <= 16'h0000;
      coeffs_in_data_log_force[5001] <= 16'h0000;
      coeffs_in_data_log_force[5002] <= 16'h0000;
      coeffs_in_data_log_force[5003] <= 16'h0000;
      coeffs_in_data_log_force[5004] <= 16'h0000;
      coeffs_in_data_log_force[5005] <= 16'h0000;
      coeffs_in_data_log_force[5006] <= 16'h0000;
      coeffs_in_data_log_force[5007] <= 16'h0000;
      coeffs_in_data_log_force[5008] <= 16'h0000;
      coeffs_in_data_log_force[5009] <= 16'h0000;
      coeffs_in_data_log_force[5010] <= 16'h0000;
      coeffs_in_data_log_force[5011] <= 16'h0000;
      coeffs_in_data_log_force[5012] <= 16'h0000;
      coeffs_in_data_log_force[5013] <= 16'h0000;
      coeffs_in_data_log_force[5014] <= 16'h0000;
      coeffs_in_data_log_force[5015] <= 16'h0000;
      coeffs_in_data_log_force[5016] <= 16'h0000;
      coeffs_in_data_log_force[5017] <= 16'h0000;
      coeffs_in_data_log_force[5018] <= 16'h0000;
      coeffs_in_data_log_force[5019] <= 16'h0000;
      coeffs_in_data_log_force[5020] <= 16'h0000;
      coeffs_in_data_log_force[5021] <= 16'h0000;
      coeffs_in_data_log_force[5022] <= 16'h0000;
      coeffs_in_data_log_force[5023] <= 16'h0000;
      coeffs_in_data_log_force[5024] <= 16'h0000;
      coeffs_in_data_log_force[5025] <= 16'h0000;
      coeffs_in_data_log_force[5026] <= 16'h0000;
      coeffs_in_data_log_force[5027] <= 16'h0000;
      coeffs_in_data_log_force[5028] <= 16'h0000;
      coeffs_in_data_log_force[5029] <= 16'h0000;
      coeffs_in_data_log_force[5030] <= 16'h0000;
      coeffs_in_data_log_force[5031] <= 16'h0000;
      coeffs_in_data_log_force[5032] <= 16'h0000;
      coeffs_in_data_log_force[5033] <= 16'h0000;
      coeffs_in_data_log_force[5034] <= 16'h0000;
      coeffs_in_data_log_force[5035] <= 16'h0000;
      coeffs_in_data_log_force[5036] <= 16'h0000;
      coeffs_in_data_log_force[5037] <= 16'h0000;
      coeffs_in_data_log_force[5038] <= 16'h0000;
      coeffs_in_data_log_force[5039] <= 16'h0000;
      coeffs_in_data_log_force[5040] <= 16'h0000;
      coeffs_in_data_log_force[5041] <= 16'h0000;
      coeffs_in_data_log_force[5042] <= 16'h0000;
      coeffs_in_data_log_force[5043] <= 16'h0000;
      coeffs_in_data_log_force[5044] <= 16'h0000;
      coeffs_in_data_log_force[5045] <= 16'h0000;
      coeffs_in_data_log_force[5046] <= 16'h0000;
      coeffs_in_data_log_force[5047] <= 16'h0000;
      coeffs_in_data_log_force[5048] <= 16'h0000;
      coeffs_in_data_log_force[5049] <= 16'h0000;
      coeffs_in_data_log_force[5050] <= 16'h0000;
      coeffs_in_data_log_force[5051] <= 16'h0000;
      coeffs_in_data_log_force[5052] <= 16'h0000;
      coeffs_in_data_log_force[5053] <= 16'h0000;
      coeffs_in_data_log_force[5054] <= 16'h0000;
      coeffs_in_data_log_force[5055] <= 16'h0000;
      coeffs_in_data_log_force[5056] <= 16'h0000;
      coeffs_in_data_log_force[5057] <= 16'h0000;
      coeffs_in_data_log_force[5058] <= 16'h0000;
      coeffs_in_data_log_force[5059] <= 16'h0000;
      coeffs_in_data_log_force[5060] <= 16'h0000;
      coeffs_in_data_log_force[5061] <= 16'h0000;
      coeffs_in_data_log_force[5062] <= 16'h0000;
      coeffs_in_data_log_force[5063] <= 16'h0000;
      coeffs_in_data_log_force[5064] <= 16'h0000;
      coeffs_in_data_log_force[5065] <= 16'h0000;
      coeffs_in_data_log_force[5066] <= 16'h0000;
      coeffs_in_data_log_force[5067] <= 16'h0000;
      coeffs_in_data_log_force[5068] <= 16'h0000;
      coeffs_in_data_log_force[5069] <= 16'h0000;
      coeffs_in_data_log_force[5070] <= 16'h0000;
      coeffs_in_data_log_force[5071] <= 16'h0000;
      coeffs_in_data_log_force[5072] <= 16'h0000;
      coeffs_in_data_log_force[5073] <= 16'h0000;
      coeffs_in_data_log_force[5074] <= 16'h0000;
      coeffs_in_data_log_force[5075] <= 16'h0000;
      coeffs_in_data_log_force[5076] <= 16'h0000;
      coeffs_in_data_log_force[5077] <= 16'h0000;
      coeffs_in_data_log_force[5078] <= 16'h0000;
      coeffs_in_data_log_force[5079] <= 16'h0000;
      coeffs_in_data_log_force[5080] <= 16'h0000;
      coeffs_in_data_log_force[5081] <= 16'h0000;
      coeffs_in_data_log_force[5082] <= 16'h0000;
      coeffs_in_data_log_force[5083] <= 16'h0000;
      coeffs_in_data_log_force[5084] <= 16'h0000;
      coeffs_in_data_log_force[5085] <= 16'h0000;
      coeffs_in_data_log_force[5086] <= 16'h0000;
      coeffs_in_data_log_force[5087] <= 16'h0000;
      coeffs_in_data_log_force[5088] <= 16'h0000;
      coeffs_in_data_log_force[5089] <= 16'h0000;
      coeffs_in_data_log_force[5090] <= 16'h0000;
      coeffs_in_data_log_force[5091] <= 16'h0000;
      coeffs_in_data_log_force[5092] <= 16'h0000;
      coeffs_in_data_log_force[5093] <= 16'h0000;
      coeffs_in_data_log_force[5094] <= 16'h0000;
      coeffs_in_data_log_force[5095] <= 16'h0000;
      coeffs_in_data_log_force[5096] <= 16'h0000;
      coeffs_in_data_log_force[5097] <= 16'h0000;
      coeffs_in_data_log_force[5098] <= 16'h0000;
      coeffs_in_data_log_force[5099] <= 16'h0000;
      coeffs_in_data_log_force[5100] <= 16'h0000;
      coeffs_in_data_log_force[5101] <= 16'h0000;
      coeffs_in_data_log_force[5102] <= 16'h0000;
      coeffs_in_data_log_force[5103] <= 16'h0000;
      coeffs_in_data_log_force[5104] <= 16'h0000;
      coeffs_in_data_log_force[5105] <= 16'h0000;
      coeffs_in_data_log_force[5106] <= 16'h0000;
      coeffs_in_data_log_force[5107] <= 16'h0000;
      coeffs_in_data_log_force[5108] <= 16'h0000;
      coeffs_in_data_log_force[5109] <= 16'h0000;
      coeffs_in_data_log_force[5110] <= 16'h0000;
      coeffs_in_data_log_force[5111] <= 16'h0000;
      coeffs_in_data_log_force[5112] <= 16'h0000;
      coeffs_in_data_log_force[5113] <= 16'h0000;
      coeffs_in_data_log_force[5114] <= 16'h0000;
      coeffs_in_data_log_force[5115] <= 16'h0000;
      coeffs_in_data_log_force[5116] <= 16'h0000;
      coeffs_in_data_log_force[5117] <= 16'h0000;
      coeffs_in_data_log_force[5118] <= 16'h0000;
      coeffs_in_data_log_force[5119] <= 16'h0000;
      coeffs_in_data_log_force[5120] <= 16'h0000;
      coeffs_in_data_log_force[5121] <= 16'h0000;
      coeffs_in_data_log_force[5122] <= 16'h0000;
      coeffs_in_data_log_force[5123] <= 16'h0000;
      coeffs_in_data_log_force[5124] <= 16'h0000;
      coeffs_in_data_log_force[5125] <= 16'h0000;
      coeffs_in_data_log_force[5126] <= 16'h0000;
      coeffs_in_data_log_force[5127] <= 16'h0000;
      coeffs_in_data_log_force[5128] <= 16'h0000;
      coeffs_in_data_log_force[5129] <= 16'h0000;
      coeffs_in_data_log_force[5130] <= 16'h0000;
      coeffs_in_data_log_force[5131] <= 16'h0000;
      coeffs_in_data_log_force[5132] <= 16'h0000;
      coeffs_in_data_log_force[5133] <= 16'h0000;
      coeffs_in_data_log_force[5134] <= 16'h0000;
      coeffs_in_data_log_force[5135] <= 16'h0000;
      coeffs_in_data_log_force[5136] <= 16'h0000;
      coeffs_in_data_log_force[5137] <= 16'h0000;
      coeffs_in_data_log_force[5138] <= 16'h0000;
      coeffs_in_data_log_force[5139] <= 16'h0000;
      coeffs_in_data_log_force[5140] <= 16'h0000;
      coeffs_in_data_log_force[5141] <= 16'h0000;
      coeffs_in_data_log_force[5142] <= 16'h0000;
      coeffs_in_data_log_force[5143] <= 16'h0000;
      coeffs_in_data_log_force[5144] <= 16'h0000;
      coeffs_in_data_log_force[5145] <= 16'h0000;
      coeffs_in_data_log_force[5146] <= 16'h0000;
      coeffs_in_data_log_force[5147] <= 16'h0000;
      coeffs_in_data_log_force[5148] <= 16'h0000;
      coeffs_in_data_log_force[5149] <= 16'h0000;
      coeffs_in_data_log_force[5150] <= 16'h0000;
      coeffs_in_data_log_force[5151] <= 16'h0000;
      coeffs_in_data_log_force[5152] <= 16'h0000;
      coeffs_in_data_log_force[5153] <= 16'h0000;
      coeffs_in_data_log_force[5154] <= 16'h0000;
      coeffs_in_data_log_force[5155] <= 16'h0000;
      coeffs_in_data_log_force[5156] <= 16'h0000;
      coeffs_in_data_log_force[5157] <= 16'h0000;
      coeffs_in_data_log_force[5158] <= 16'h0000;
      coeffs_in_data_log_force[5159] <= 16'h0000;
      coeffs_in_data_log_force[5160] <= 16'h0000;
      coeffs_in_data_log_force[5161] <= 16'h0000;
      coeffs_in_data_log_force[5162] <= 16'h0000;
      coeffs_in_data_log_force[5163] <= 16'h0000;
      coeffs_in_data_log_force[5164] <= 16'h0000;
      coeffs_in_data_log_force[5165] <= 16'h0000;
      coeffs_in_data_log_force[5166] <= 16'h0000;
      coeffs_in_data_log_force[5167] <= 16'h0000;
      coeffs_in_data_log_force[5168] <= 16'h0000;
      coeffs_in_data_log_force[5169] <= 16'h0000;
      coeffs_in_data_log_force[5170] <= 16'h0000;
      coeffs_in_data_log_force[5171] <= 16'h0000;
      coeffs_in_data_log_force[5172] <= 16'h0000;
      coeffs_in_data_log_force[5173] <= 16'h0000;
      coeffs_in_data_log_force[5174] <= 16'h0000;
      coeffs_in_data_log_force[5175] <= 16'h0000;
      coeffs_in_data_log_force[5176] <= 16'h0000;
      coeffs_in_data_log_force[5177] <= 16'h0000;
      coeffs_in_data_log_force[5178] <= 16'h0000;
      coeffs_in_data_log_force[5179] <= 16'h0000;
      coeffs_in_data_log_force[5180] <= 16'h0000;
      coeffs_in_data_log_force[5181] <= 16'h0000;
      coeffs_in_data_log_force[5182] <= 16'h0000;
      coeffs_in_data_log_force[5183] <= 16'h0000;
      coeffs_in_data_log_force[5184] <= 16'h0000;
      coeffs_in_data_log_force[5185] <= 16'h0000;
      coeffs_in_data_log_force[5186] <= 16'h0000;
      coeffs_in_data_log_force[5187] <= 16'h0000;
      coeffs_in_data_log_force[5188] <= 16'h0000;
      coeffs_in_data_log_force[5189] <= 16'h0000;
      coeffs_in_data_log_force[5190] <= 16'h0000;
      coeffs_in_data_log_force[5191] <= 16'h0000;
      coeffs_in_data_log_force[5192] <= 16'h0000;
      coeffs_in_data_log_force[5193] <= 16'h0000;
      coeffs_in_data_log_force[5194] <= 16'h0000;
      coeffs_in_data_log_force[5195] <= 16'h0000;
      coeffs_in_data_log_force[5196] <= 16'h0000;
      coeffs_in_data_log_force[5197] <= 16'h0000;
      coeffs_in_data_log_force[5198] <= 16'h0000;
      coeffs_in_data_log_force[5199] <= 16'h0000;
      coeffs_in_data_log_force[5200] <= 16'h0000;
      coeffs_in_data_log_force[5201] <= 16'h0000;
      coeffs_in_data_log_force[5202] <= 16'h0000;
      coeffs_in_data_log_force[5203] <= 16'h0000;
      coeffs_in_data_log_force[5204] <= 16'h0000;
      coeffs_in_data_log_force[5205] <= 16'h0000;
      coeffs_in_data_log_force[5206] <= 16'h0000;
      coeffs_in_data_log_force[5207] <= 16'h0000;
      coeffs_in_data_log_force[5208] <= 16'h0000;
      coeffs_in_data_log_force[5209] <= 16'h0000;
      coeffs_in_data_log_force[5210] <= 16'h0000;
      coeffs_in_data_log_force[5211] <= 16'h0000;
      coeffs_in_data_log_force[5212] <= 16'h0000;
      coeffs_in_data_log_force[5213] <= 16'h0000;
      coeffs_in_data_log_force[5214] <= 16'h0000;
      coeffs_in_data_log_force[5215] <= 16'h0000;
      coeffs_in_data_log_force[5216] <= 16'h0000;
      coeffs_in_data_log_force[5217] <= 16'h0000;
      coeffs_in_data_log_force[5218] <= 16'h0000;
      coeffs_in_data_log_force[5219] <= 16'h0000;
      coeffs_in_data_log_force[5220] <= 16'h0000;
      coeffs_in_data_log_force[5221] <= 16'h0000;
      coeffs_in_data_log_force[5222] <= 16'h0000;
      coeffs_in_data_log_force[5223] <= 16'h0000;
      coeffs_in_data_log_force[5224] <= 16'h0000;
      coeffs_in_data_log_force[5225] <= 16'h0000;
      coeffs_in_data_log_force[5226] <= 16'h0000;
      coeffs_in_data_log_force[5227] <= 16'h0000;
      coeffs_in_data_log_force[5228] <= 16'h0000;
      coeffs_in_data_log_force[5229] <= 16'h0000;
      coeffs_in_data_log_force[5230] <= 16'h0000;
      coeffs_in_data_log_force[5231] <= 16'h0000;
      coeffs_in_data_log_force[5232] <= 16'h0000;
      coeffs_in_data_log_force[5233] <= 16'h0000;
      coeffs_in_data_log_force[5234] <= 16'h0000;
      coeffs_in_data_log_force[5235] <= 16'h0000;
      coeffs_in_data_log_force[5236] <= 16'h0000;
      coeffs_in_data_log_force[5237] <= 16'h0000;
      coeffs_in_data_log_force[5238] <= 16'h0000;
      coeffs_in_data_log_force[5239] <= 16'h0000;
      coeffs_in_data_log_force[5240] <= 16'h0000;
      coeffs_in_data_log_force[5241] <= 16'h0000;
      coeffs_in_data_log_force[5242] <= 16'h0000;
      coeffs_in_data_log_force[5243] <= 16'h0000;
      coeffs_in_data_log_force[5244] <= 16'h0000;
      coeffs_in_data_log_force[5245] <= 16'h0000;
      coeffs_in_data_log_force[5246] <= 16'h0000;
      coeffs_in_data_log_force[5247] <= 16'h0000;
      coeffs_in_data_log_force[5248] <= 16'h0000;
      coeffs_in_data_log_force[5249] <= 16'h0000;
      coeffs_in_data_log_force[5250] <= 16'h0000;
      coeffs_in_data_log_force[5251] <= 16'h0000;
      coeffs_in_data_log_force[5252] <= 16'h0000;
      coeffs_in_data_log_force[5253] <= 16'h0000;
      coeffs_in_data_log_force[5254] <= 16'h0000;
      coeffs_in_data_log_force[5255] <= 16'h0000;
      coeffs_in_data_log_force[5256] <= 16'h0000;
      coeffs_in_data_log_force[5257] <= 16'h0000;
      coeffs_in_data_log_force[5258] <= 16'h0000;
      coeffs_in_data_log_force[5259] <= 16'h0000;
      coeffs_in_data_log_force[5260] <= 16'h0000;
      coeffs_in_data_log_force[5261] <= 16'h0000;
      coeffs_in_data_log_force[5262] <= 16'h0000;
      coeffs_in_data_log_force[5263] <= 16'h0000;
      coeffs_in_data_log_force[5264] <= 16'h0000;
      coeffs_in_data_log_force[5265] <= 16'h0000;
      coeffs_in_data_log_force[5266] <= 16'h0000;
      coeffs_in_data_log_force[5267] <= 16'h0000;
      coeffs_in_data_log_force[5268] <= 16'h0000;
      coeffs_in_data_log_force[5269] <= 16'h0000;
      coeffs_in_data_log_force[5270] <= 16'h0000;
      coeffs_in_data_log_force[5271] <= 16'h0000;
      coeffs_in_data_log_force[5272] <= 16'h0000;
      coeffs_in_data_log_force[5273] <= 16'h0000;
      coeffs_in_data_log_force[5274] <= 16'h0000;
      coeffs_in_data_log_force[5275] <= 16'h0000;
      coeffs_in_data_log_force[5276] <= 16'h0000;
      coeffs_in_data_log_force[5277] <= 16'h0000;
      coeffs_in_data_log_force[5278] <= 16'h0000;
      coeffs_in_data_log_force[5279] <= 16'h0000;
      coeffs_in_data_log_force[5280] <= 16'h0000;
      coeffs_in_data_log_force[5281] <= 16'h0000;
      coeffs_in_data_log_force[5282] <= 16'h0000;
      coeffs_in_data_log_force[5283] <= 16'h0000;
      coeffs_in_data_log_force[5284] <= 16'h0000;
      coeffs_in_data_log_force[5285] <= 16'h0000;
      coeffs_in_data_log_force[5286] <= 16'h0000;
      coeffs_in_data_log_force[5287] <= 16'h0000;
      coeffs_in_data_log_force[5288] <= 16'h0000;
      coeffs_in_data_log_force[5289] <= 16'h0000;
      coeffs_in_data_log_force[5290] <= 16'h0000;
      coeffs_in_data_log_force[5291] <= 16'h0000;
      coeffs_in_data_log_force[5292] <= 16'h0000;
      coeffs_in_data_log_force[5293] <= 16'h0000;
      coeffs_in_data_log_force[5294] <= 16'h0000;
      coeffs_in_data_log_force[5295] <= 16'h0000;
      coeffs_in_data_log_force[5296] <= 16'h0000;
      coeffs_in_data_log_force[5297] <= 16'h0000;
      coeffs_in_data_log_force[5298] <= 16'h0000;
      coeffs_in_data_log_force[5299] <= 16'h0000;
      coeffs_in_data_log_force[5300] <= 16'h0000;
      coeffs_in_data_log_force[5301] <= 16'h0000;
      coeffs_in_data_log_force[5302] <= 16'h0000;
      coeffs_in_data_log_force[5303] <= 16'h0000;
      coeffs_in_data_log_force[5304] <= 16'h0000;
      coeffs_in_data_log_force[5305] <= 16'h0000;
      coeffs_in_data_log_force[5306] <= 16'h0000;
      coeffs_in_data_log_force[5307] <= 16'h0000;
      coeffs_in_data_log_force[5308] <= 16'h0000;
      coeffs_in_data_log_force[5309] <= 16'h0000;
      coeffs_in_data_log_force[5310] <= 16'h0000;
      coeffs_in_data_log_force[5311] <= 16'h0000;
      coeffs_in_data_log_force[5312] <= 16'h0000;
      coeffs_in_data_log_force[5313] <= 16'h0000;
      coeffs_in_data_log_force[5314] <= 16'h0000;
      coeffs_in_data_log_force[5315] <= 16'h0000;
      coeffs_in_data_log_force[5316] <= 16'h0000;
      coeffs_in_data_log_force[5317] <= 16'h0000;
      coeffs_in_data_log_force[5318] <= 16'h0000;
      coeffs_in_data_log_force[5319] <= 16'h0000;
      coeffs_in_data_log_force[5320] <= 16'h0000;
      coeffs_in_data_log_force[5321] <= 16'h0000;
      coeffs_in_data_log_force[5322] <= 16'h0000;
      coeffs_in_data_log_force[5323] <= 16'h0000;
      coeffs_in_data_log_force[5324] <= 16'h0000;
      coeffs_in_data_log_force[5325] <= 16'h0000;
      coeffs_in_data_log_force[5326] <= 16'h0000;
      coeffs_in_data_log_force[5327] <= 16'h0000;
      coeffs_in_data_log_force[5328] <= 16'h0000;
      coeffs_in_data_log_force[5329] <= 16'h0000;
      coeffs_in_data_log_force[5330] <= 16'h0000;
      coeffs_in_data_log_force[5331] <= 16'h0000;
      coeffs_in_data_log_force[5332] <= 16'h0000;
      coeffs_in_data_log_force[5333] <= 16'h0000;
      coeffs_in_data_log_force[5334] <= 16'h0000;
      coeffs_in_data_log_force[5335] <= 16'h0000;
      coeffs_in_data_log_force[5336] <= 16'h0000;
      coeffs_in_data_log_force[5337] <= 16'h0000;
      coeffs_in_data_log_force[5338] <= 16'h0000;
      coeffs_in_data_log_force[5339] <= 16'h0000;
      coeffs_in_data_log_force[5340] <= 16'h0000;
      coeffs_in_data_log_force[5341] <= 16'h0000;
      coeffs_in_data_log_force[5342] <= 16'h0000;
      coeffs_in_data_log_force[5343] <= 16'h0000;
      coeffs_in_data_log_force[5344] <= 16'h0000;
      coeffs_in_data_log_force[5345] <= 16'h0000;
      coeffs_in_data_log_force[5346] <= 16'h0000;
      coeffs_in_data_log_force[5347] <= 16'h0000;
      coeffs_in_data_log_force[5348] <= 16'h0000;
      coeffs_in_data_log_force[5349] <= 16'h0000;
      coeffs_in_data_log_force[5350] <= 16'h0000;
      coeffs_in_data_log_force[5351] <= 16'h0000;
      coeffs_in_data_log_force[5352] <= 16'h0000;
      coeffs_in_data_log_force[5353] <= 16'h0000;
      coeffs_in_data_log_force[5354] <= 16'h0000;
      coeffs_in_data_log_force[5355] <= 16'h0000;
      coeffs_in_data_log_force[5356] <= 16'h0000;
      coeffs_in_data_log_force[5357] <= 16'h0000;
      coeffs_in_data_log_force[5358] <= 16'h0000;
      coeffs_in_data_log_force[5359] <= 16'h0000;
      coeffs_in_data_log_force[5360] <= 16'h0000;
      coeffs_in_data_log_force[5361] <= 16'h0000;
      coeffs_in_data_log_force[5362] <= 16'h0000;
      coeffs_in_data_log_force[5363] <= 16'h0000;
      coeffs_in_data_log_force[5364] <= 16'h0000;
      coeffs_in_data_log_force[5365] <= 16'h0000;
      coeffs_in_data_log_force[5366] <= 16'h0000;
      coeffs_in_data_log_force[5367] <= 16'h0000;
      coeffs_in_data_log_force[5368] <= 16'h0000;
      coeffs_in_data_log_force[5369] <= 16'h0000;
      coeffs_in_data_log_force[5370] <= 16'h0000;
      coeffs_in_data_log_force[5371] <= 16'h0000;
      coeffs_in_data_log_force[5372] <= 16'h0000;
      coeffs_in_data_log_force[5373] <= 16'h0000;
      coeffs_in_data_log_force[5374] <= 16'h0000;
      coeffs_in_data_log_force[5375] <= 16'h0000;
      coeffs_in_data_log_force[5376] <= 16'h0000;
      coeffs_in_data_log_force[5377] <= 16'h0000;
      coeffs_in_data_log_force[5378] <= 16'h0000;
      coeffs_in_data_log_force[5379] <= 16'h0000;
      coeffs_in_data_log_force[5380] <= 16'h0000;
      coeffs_in_data_log_force[5381] <= 16'h0000;
      coeffs_in_data_log_force[5382] <= 16'h0000;
      coeffs_in_data_log_force[5383] <= 16'h0000;
      coeffs_in_data_log_force[5384] <= 16'h0000;
      coeffs_in_data_log_force[5385] <= 16'h0000;
      coeffs_in_data_log_force[5386] <= 16'h0000;
      coeffs_in_data_log_force[5387] <= 16'h0000;
      coeffs_in_data_log_force[5388] <= 16'h0000;
      coeffs_in_data_log_force[5389] <= 16'h0000;
      coeffs_in_data_log_force[5390] <= 16'h0000;
      coeffs_in_data_log_force[5391] <= 16'h0000;
      coeffs_in_data_log_force[5392] <= 16'h0000;
      coeffs_in_data_log_force[5393] <= 16'h0000;
      coeffs_in_data_log_force[5394] <= 16'h0000;
      coeffs_in_data_log_force[5395] <= 16'h0000;
      coeffs_in_data_log_force[5396] <= 16'h0000;
      coeffs_in_data_log_force[5397] <= 16'h0000;
      coeffs_in_data_log_force[5398] <= 16'h0000;
      coeffs_in_data_log_force[5399] <= 16'h0000;
      coeffs_in_data_log_force[5400] <= 16'h0000;
      coeffs_in_data_log_force[5401] <= 16'h0000;
      coeffs_in_data_log_force[5402] <= 16'h0000;
      coeffs_in_data_log_force[5403] <= 16'h0000;
      coeffs_in_data_log_force[5404] <= 16'h0000;
      coeffs_in_data_log_force[5405] <= 16'h0000;
      coeffs_in_data_log_force[5406] <= 16'h0000;
      coeffs_in_data_log_force[5407] <= 16'h0000;
      coeffs_in_data_log_force[5408] <= 16'h0000;
      coeffs_in_data_log_force[5409] <= 16'h0000;
      coeffs_in_data_log_force[5410] <= 16'h0000;
      coeffs_in_data_log_force[5411] <= 16'h0000;
      coeffs_in_data_log_force[5412] <= 16'h0000;
      coeffs_in_data_log_force[5413] <= 16'h0000;
      coeffs_in_data_log_force[5414] <= 16'h0000;
      coeffs_in_data_log_force[5415] <= 16'h0000;
      coeffs_in_data_log_force[5416] <= 16'h0000;
      coeffs_in_data_log_force[5417] <= 16'h0000;
      coeffs_in_data_log_force[5418] <= 16'h0000;
      coeffs_in_data_log_force[5419] <= 16'h0000;
      coeffs_in_data_log_force[5420] <= 16'h0000;
      coeffs_in_data_log_force[5421] <= 16'h0000;
      coeffs_in_data_log_force[5422] <= 16'h0000;
      coeffs_in_data_log_force[5423] <= 16'h0000;
      coeffs_in_data_log_force[5424] <= 16'h0000;
      coeffs_in_data_log_force[5425] <= 16'h0000;
      coeffs_in_data_log_force[5426] <= 16'h0000;
      coeffs_in_data_log_force[5427] <= 16'h0000;
      coeffs_in_data_log_force[5428] <= 16'h0000;
      coeffs_in_data_log_force[5429] <= 16'h0000;
      coeffs_in_data_log_force[5430] <= 16'h0000;
      coeffs_in_data_log_force[5431] <= 16'h0000;
      coeffs_in_data_log_force[5432] <= 16'h0000;
      coeffs_in_data_log_force[5433] <= 16'h0000;
      coeffs_in_data_log_force[5434] <= 16'h0000;
      coeffs_in_data_log_force[5435] <= 16'h0000;
      coeffs_in_data_log_force[5436] <= 16'h0000;
      coeffs_in_data_log_force[5437] <= 16'h0000;
      coeffs_in_data_log_force[5438] <= 16'h0000;
      coeffs_in_data_log_force[5439] <= 16'h0000;
      coeffs_in_data_log_force[5440] <= 16'h0000;
      coeffs_in_data_log_force[5441] <= 16'h0000;
      coeffs_in_data_log_force[5442] <= 16'h0000;
      coeffs_in_data_log_force[5443] <= 16'h0000;
      coeffs_in_data_log_force[5444] <= 16'h0000;
      coeffs_in_data_log_force[5445] <= 16'h0000;
      coeffs_in_data_log_force[5446] <= 16'h0000;
      coeffs_in_data_log_force[5447] <= 16'h0000;
      coeffs_in_data_log_force[5448] <= 16'h0000;
      coeffs_in_data_log_force[5449] <= 16'h0000;
      coeffs_in_data_log_force[5450] <= 16'h0000;
      coeffs_in_data_log_force[5451] <= 16'h0000;
      coeffs_in_data_log_force[5452] <= 16'h0000;
      coeffs_in_data_log_force[5453] <= 16'h0000;
      coeffs_in_data_log_force[5454] <= 16'h0000;
      coeffs_in_data_log_force[5455] <= 16'h0000;
      coeffs_in_data_log_force[5456] <= 16'h0000;
      coeffs_in_data_log_force[5457] <= 16'h0000;
      coeffs_in_data_log_force[5458] <= 16'h0000;
      coeffs_in_data_log_force[5459] <= 16'h0000;
      coeffs_in_data_log_force[5460] <= 16'h0000;
      coeffs_in_data_log_force[5461] <= 16'h0000;
      coeffs_in_data_log_force[5462] <= 16'h0000;
      coeffs_in_data_log_force[5463] <= 16'h0000;
      coeffs_in_data_log_force[5464] <= 16'h0000;
      coeffs_in_data_log_force[5465] <= 16'h0000;
      coeffs_in_data_log_force[5466] <= 16'h0000;
      coeffs_in_data_log_force[5467] <= 16'h0000;
      coeffs_in_data_log_force[5468] <= 16'h0000;
      coeffs_in_data_log_force[5469] <= 16'h0000;
      coeffs_in_data_log_force[5470] <= 16'h0000;
      coeffs_in_data_log_force[5471] <= 16'h0000;
      coeffs_in_data_log_force[5472] <= 16'h0000;
      coeffs_in_data_log_force[5473] <= 16'h0000;
      coeffs_in_data_log_force[5474] <= 16'h0000;
      coeffs_in_data_log_force[5475] <= 16'h0000;
      coeffs_in_data_log_force[5476] <= 16'h0000;
      coeffs_in_data_log_force[5477] <= 16'h0000;
      coeffs_in_data_log_force[5478] <= 16'h0000;
      coeffs_in_data_log_force[5479] <= 16'h0000;
      coeffs_in_data_log_force[5480] <= 16'h0000;
      coeffs_in_data_log_force[5481] <= 16'h0000;
      coeffs_in_data_log_force[5482] <= 16'h0000;
      coeffs_in_data_log_force[5483] <= 16'h0000;
      coeffs_in_data_log_force[5484] <= 16'h0000;
      coeffs_in_data_log_force[5485] <= 16'h0000;
      coeffs_in_data_log_force[5486] <= 16'h0000;
      coeffs_in_data_log_force[5487] <= 16'h0000;
      coeffs_in_data_log_force[5488] <= 16'h0000;
      coeffs_in_data_log_force[5489] <= 16'h0000;
      coeffs_in_data_log_force[5490] <= 16'h0000;
      coeffs_in_data_log_force[5491] <= 16'h0000;
      coeffs_in_data_log_force[5492] <= 16'h0000;
      coeffs_in_data_log_force[5493] <= 16'h0000;
      coeffs_in_data_log_force[5494] <= 16'h0000;
      coeffs_in_data_log_force[5495] <= 16'h0000;
      coeffs_in_data_log_force[5496] <= 16'h0000;
      coeffs_in_data_log_force[5497] <= 16'h0000;
      coeffs_in_data_log_force[5498] <= 16'h0000;
      coeffs_in_data_log_force[5499] <= 16'h0000;
      coeffs_in_data_log_force[5500] <= 16'h0000;
      coeffs_in_data_log_force[5501] <= 16'h0000;
      coeffs_in_data_log_force[5502] <= 16'h0000;
      coeffs_in_data_log_force[5503] <= 16'h0000;
      coeffs_in_data_log_force[5504] <= 16'h0000;
      coeffs_in_data_log_force[5505] <= 16'h0000;
      coeffs_in_data_log_force[5506] <= 16'h0000;
      coeffs_in_data_log_force[5507] <= 16'h0000;
      coeffs_in_data_log_force[5508] <= 16'h0000;
      coeffs_in_data_log_force[5509] <= 16'h0000;
      coeffs_in_data_log_force[5510] <= 16'h0000;
      coeffs_in_data_log_force[5511] <= 16'h0000;
      coeffs_in_data_log_force[5512] <= 16'h0000;
      coeffs_in_data_log_force[5513] <= 16'h0000;
      coeffs_in_data_log_force[5514] <= 16'h0000;
      coeffs_in_data_log_force[5515] <= 16'h0000;
      coeffs_in_data_log_force[5516] <= 16'h0000;
      coeffs_in_data_log_force[5517] <= 16'h0000;
      coeffs_in_data_log_force[5518] <= 16'h0000;
      coeffs_in_data_log_force[5519] <= 16'h0000;
      coeffs_in_data_log_force[5520] <= 16'h0000;
      coeffs_in_data_log_force[5521] <= 16'h0000;
      coeffs_in_data_log_force[5522] <= 16'h0000;
      coeffs_in_data_log_force[5523] <= 16'h0000;
      coeffs_in_data_log_force[5524] <= 16'h0000;
      coeffs_in_data_log_force[5525] <= 16'h0000;
      coeffs_in_data_log_force[5526] <= 16'h0000;
      coeffs_in_data_log_force[5527] <= 16'h0000;
      coeffs_in_data_log_force[5528] <= 16'h0000;
      coeffs_in_data_log_force[5529] <= 16'h0000;
      coeffs_in_data_log_force[5530] <= 16'h0000;
      coeffs_in_data_log_force[5531] <= 16'h0000;
      coeffs_in_data_log_force[5532] <= 16'h0000;
      coeffs_in_data_log_force[5533] <= 16'h0000;
      coeffs_in_data_log_force[5534] <= 16'h0000;
      coeffs_in_data_log_force[5535] <= 16'h0000;
      coeffs_in_data_log_force[5536] <= 16'h0000;
      coeffs_in_data_log_force[5537] <= 16'h0000;
      coeffs_in_data_log_force[5538] <= 16'h0000;
      coeffs_in_data_log_force[5539] <= 16'h0000;
      coeffs_in_data_log_force[5540] <= 16'h0000;
      coeffs_in_data_log_force[5541] <= 16'h0000;
      coeffs_in_data_log_force[5542] <= 16'h0000;
      coeffs_in_data_log_force[5543] <= 16'h0000;
      coeffs_in_data_log_force[5544] <= 16'h0000;
      coeffs_in_data_log_force[5545] <= 16'h0000;
      coeffs_in_data_log_force[5546] <= 16'h0000;
      coeffs_in_data_log_force[5547] <= 16'h0000;
      coeffs_in_data_log_force[5548] <= 16'h0000;
      coeffs_in_data_log_force[5549] <= 16'h0000;
      coeffs_in_data_log_force[5550] <= 16'h0000;
      coeffs_in_data_log_force[5551] <= 16'h0000;
      coeffs_in_data_log_force[5552] <= 16'h0000;
      coeffs_in_data_log_force[5553] <= 16'h0000;
      coeffs_in_data_log_force[5554] <= 16'h0000;
      coeffs_in_data_log_force[5555] <= 16'h0000;
      coeffs_in_data_log_force[5556] <= 16'h0000;
      coeffs_in_data_log_force[5557] <= 16'h0000;
      coeffs_in_data_log_force[5558] <= 16'h0000;
      coeffs_in_data_log_force[5559] <= 16'h0000;
      coeffs_in_data_log_force[5560] <= 16'h0000;
      coeffs_in_data_log_force[5561] <= 16'h0000;
      coeffs_in_data_log_force[5562] <= 16'h0000;
      coeffs_in_data_log_force[5563] <= 16'h0000;
      coeffs_in_data_log_force[5564] <= 16'h0000;
      coeffs_in_data_log_force[5565] <= 16'h0000;
      coeffs_in_data_log_force[5566] <= 16'h0000;
      coeffs_in_data_log_force[5567] <= 16'h0000;
      coeffs_in_data_log_force[5568] <= 16'h0000;
      coeffs_in_data_log_force[5569] <= 16'h0000;
      coeffs_in_data_log_force[5570] <= 16'h0000;
      coeffs_in_data_log_force[5571] <= 16'h0000;
      coeffs_in_data_log_force[5572] <= 16'h0000;
      coeffs_in_data_log_force[5573] <= 16'h0000;
      coeffs_in_data_log_force[5574] <= 16'h0000;
      coeffs_in_data_log_force[5575] <= 16'h0000;
      coeffs_in_data_log_force[5576] <= 16'h0000;
      coeffs_in_data_log_force[5577] <= 16'h0000;
      coeffs_in_data_log_force[5578] <= 16'h0000;
      coeffs_in_data_log_force[5579] <= 16'h0000;
      coeffs_in_data_log_force[5580] <= 16'h0000;
      coeffs_in_data_log_force[5581] <= 16'h0000;
      coeffs_in_data_log_force[5582] <= 16'h0000;
      coeffs_in_data_log_force[5583] <= 16'h0000;
      coeffs_in_data_log_force[5584] <= 16'h0000;
      coeffs_in_data_log_force[5585] <= 16'h0000;
      coeffs_in_data_log_force[5586] <= 16'h0000;
      coeffs_in_data_log_force[5587] <= 16'h0000;
      coeffs_in_data_log_force[5588] <= 16'h0000;
      coeffs_in_data_log_force[5589] <= 16'h0000;
      coeffs_in_data_log_force[5590] <= 16'h0000;
      coeffs_in_data_log_force[5591] <= 16'h0000;
      coeffs_in_data_log_force[5592] <= 16'h0000;
      coeffs_in_data_log_force[5593] <= 16'h0000;
      coeffs_in_data_log_force[5594] <= 16'h0000;
      coeffs_in_data_log_force[5595] <= 16'h0000;
      coeffs_in_data_log_force[5596] <= 16'h0000;
      coeffs_in_data_log_force[5597] <= 16'h0000;
      coeffs_in_data_log_force[5598] <= 16'h0000;
      coeffs_in_data_log_force[5599] <= 16'h0000;
      coeffs_in_data_log_force[5600] <= 16'h0000;
      coeffs_in_data_log_force[5601] <= 16'h0000;
      coeffs_in_data_log_force[5602] <= 16'h0000;
      coeffs_in_data_log_force[5603] <= 16'h0000;
      coeffs_in_data_log_force[5604] <= 16'h0000;
      coeffs_in_data_log_force[5605] <= 16'h0000;
      coeffs_in_data_log_force[5606] <= 16'h0000;
      coeffs_in_data_log_force[5607] <= 16'h0000;
      coeffs_in_data_log_force[5608] <= 16'h0000;
      coeffs_in_data_log_force[5609] <= 16'h0000;
      coeffs_in_data_log_force[5610] <= 16'h0000;
      coeffs_in_data_log_force[5611] <= 16'h0000;
      coeffs_in_data_log_force[5612] <= 16'h0000;
      coeffs_in_data_log_force[5613] <= 16'h0000;
      coeffs_in_data_log_force[5614] <= 16'h0000;
      coeffs_in_data_log_force[5615] <= 16'h0000;
      coeffs_in_data_log_force[5616] <= 16'h0000;
      coeffs_in_data_log_force[5617] <= 16'h0000;
      coeffs_in_data_log_force[5618] <= 16'h0000;
      coeffs_in_data_log_force[5619] <= 16'h0000;
      coeffs_in_data_log_force[5620] <= 16'h0000;
      coeffs_in_data_log_force[5621] <= 16'h0000;
      coeffs_in_data_log_force[5622] <= 16'h0000;
      coeffs_in_data_log_force[5623] <= 16'h0000;
      coeffs_in_data_log_force[5624] <= 16'h0000;
      coeffs_in_data_log_force[5625] <= 16'h0000;
      coeffs_in_data_log_force[5626] <= 16'h0000;
      coeffs_in_data_log_force[5627] <= 16'h0000;
      coeffs_in_data_log_force[5628] <= 16'h0000;
      coeffs_in_data_log_force[5629] <= 16'h0000;
      coeffs_in_data_log_force[5630] <= 16'h0000;
      coeffs_in_data_log_force[5631] <= 16'h0000;
      coeffs_in_data_log_force[5632] <= 16'h0000;
      coeffs_in_data_log_force[5633] <= 16'h0000;
      coeffs_in_data_log_force[5634] <= 16'h0000;
      coeffs_in_data_log_force[5635] <= 16'h0000;
      coeffs_in_data_log_force[5636] <= 16'h0000;
      coeffs_in_data_log_force[5637] <= 16'h0000;
      coeffs_in_data_log_force[5638] <= 16'h0000;
      coeffs_in_data_log_force[5639] <= 16'h0000;
      coeffs_in_data_log_force[5640] <= 16'h0000;
      coeffs_in_data_log_force[5641] <= 16'h0000;
      coeffs_in_data_log_force[5642] <= 16'h0000;
      coeffs_in_data_log_force[5643] <= 16'h0000;
      coeffs_in_data_log_force[5644] <= 16'h0000;
      coeffs_in_data_log_force[5645] <= 16'h0000;
      coeffs_in_data_log_force[5646] <= 16'h0000;
      coeffs_in_data_log_force[5647] <= 16'h0000;
      coeffs_in_data_log_force[5648] <= 16'h0000;
      coeffs_in_data_log_force[5649] <= 16'h0000;
      coeffs_in_data_log_force[5650] <= 16'h0000;
      coeffs_in_data_log_force[5651] <= 16'h0000;
      coeffs_in_data_log_force[5652] <= 16'h0000;
      coeffs_in_data_log_force[5653] <= 16'h0000;
      coeffs_in_data_log_force[5654] <= 16'h0000;
      coeffs_in_data_log_force[5655] <= 16'h0000;
      coeffs_in_data_log_force[5656] <= 16'h0000;
      coeffs_in_data_log_force[5657] <= 16'h0000;
      coeffs_in_data_log_force[5658] <= 16'h0000;
      coeffs_in_data_log_force[5659] <= 16'h0000;
      coeffs_in_data_log_force[5660] <= 16'h0000;
      coeffs_in_data_log_force[5661] <= 16'h0000;
      coeffs_in_data_log_force[5662] <= 16'h0000;
      coeffs_in_data_log_force[5663] <= 16'h0000;
      coeffs_in_data_log_force[5664] <= 16'h0000;
      coeffs_in_data_log_force[5665] <= 16'h0000;
      coeffs_in_data_log_force[5666] <= 16'h0000;
      coeffs_in_data_log_force[5667] <= 16'h0000;
      coeffs_in_data_log_force[5668] <= 16'h0000;
      coeffs_in_data_log_force[5669] <= 16'h0000;
      coeffs_in_data_log_force[5670] <= 16'h0000;
      coeffs_in_data_log_force[5671] <= 16'h0000;
      coeffs_in_data_log_force[5672] <= 16'h0000;
      coeffs_in_data_log_force[5673] <= 16'h0000;
      coeffs_in_data_log_force[5674] <= 16'h0000;
      coeffs_in_data_log_force[5675] <= 16'h0000;
      coeffs_in_data_log_force[5676] <= 16'h0000;
      coeffs_in_data_log_force[5677] <= 16'h0000;
      coeffs_in_data_log_force[5678] <= 16'h0000;
      coeffs_in_data_log_force[5679] <= 16'h0000;
      coeffs_in_data_log_force[5680] <= 16'h0000;
      coeffs_in_data_log_force[5681] <= 16'h0000;
      coeffs_in_data_log_force[5682] <= 16'h0000;
      coeffs_in_data_log_force[5683] <= 16'h0000;
      coeffs_in_data_log_force[5684] <= 16'h0000;
      coeffs_in_data_log_force[5685] <= 16'h0000;
      coeffs_in_data_log_force[5686] <= 16'h0000;
      coeffs_in_data_log_force[5687] <= 16'h0000;
      coeffs_in_data_log_force[5688] <= 16'h0000;
      coeffs_in_data_log_force[5689] <= 16'h0000;
      coeffs_in_data_log_force[5690] <= 16'h0000;
      coeffs_in_data_log_force[5691] <= 16'h0000;
      coeffs_in_data_log_force[5692] <= 16'h0000;
      coeffs_in_data_log_force[5693] <= 16'h0000;
      coeffs_in_data_log_force[5694] <= 16'h0000;
      coeffs_in_data_log_force[5695] <= 16'h0000;
      coeffs_in_data_log_force[5696] <= 16'h0000;
      coeffs_in_data_log_force[5697] <= 16'h0000;
      coeffs_in_data_log_force[5698] <= 16'h0000;
      coeffs_in_data_log_force[5699] <= 16'h0000;
      coeffs_in_data_log_force[5700] <= 16'h0000;
      coeffs_in_data_log_force[5701] <= 16'h0000;
      coeffs_in_data_log_force[5702] <= 16'h0000;
      coeffs_in_data_log_force[5703] <= 16'h0000;
      coeffs_in_data_log_force[5704] <= 16'h0000;
      coeffs_in_data_log_force[5705] <= 16'h0000;
      coeffs_in_data_log_force[5706] <= 16'h0000;
      coeffs_in_data_log_force[5707] <= 16'h0000;
      coeffs_in_data_log_force[5708] <= 16'h0000;
      coeffs_in_data_log_force[5709] <= 16'h0000;
      coeffs_in_data_log_force[5710] <= 16'h0000;
      coeffs_in_data_log_force[5711] <= 16'h0000;
      coeffs_in_data_log_force[5712] <= 16'h0000;
      coeffs_in_data_log_force[5713] <= 16'h0000;
      coeffs_in_data_log_force[5714] <= 16'h0000;
      coeffs_in_data_log_force[5715] <= 16'h0000;
      coeffs_in_data_log_force[5716] <= 16'h0000;
      coeffs_in_data_log_force[5717] <= 16'h0000;
      coeffs_in_data_log_force[5718] <= 16'h0000;
      coeffs_in_data_log_force[5719] <= 16'h0000;
      coeffs_in_data_log_force[5720] <= 16'h0000;
      coeffs_in_data_log_force[5721] <= 16'h0000;
      coeffs_in_data_log_force[5722] <= 16'h0000;
      coeffs_in_data_log_force[5723] <= 16'h0000;
      coeffs_in_data_log_force[5724] <= 16'h0000;
      coeffs_in_data_log_force[5725] <= 16'h0000;
      coeffs_in_data_log_force[5726] <= 16'h0000;
      coeffs_in_data_log_force[5727] <= 16'h0000;
      coeffs_in_data_log_force[5728] <= 16'h0000;
      coeffs_in_data_log_force[5729] <= 16'h0000;
      coeffs_in_data_log_force[5730] <= 16'h0000;
      coeffs_in_data_log_force[5731] <= 16'h0000;
      coeffs_in_data_log_force[5732] <= 16'h0000;
      coeffs_in_data_log_force[5733] <= 16'h0000;
      coeffs_in_data_log_force[5734] <= 16'h0000;
      coeffs_in_data_log_force[5735] <= 16'h0000;
      coeffs_in_data_log_force[5736] <= 16'h0000;
      coeffs_in_data_log_force[5737] <= 16'h0000;
      coeffs_in_data_log_force[5738] <= 16'h0000;
      coeffs_in_data_log_force[5739] <= 16'h0000;
      coeffs_in_data_log_force[5740] <= 16'h0000;
      coeffs_in_data_log_force[5741] <= 16'h0000;
      coeffs_in_data_log_force[5742] <= 16'h0000;
      coeffs_in_data_log_force[5743] <= 16'h0000;
      coeffs_in_data_log_force[5744] <= 16'h0000;
      coeffs_in_data_log_force[5745] <= 16'h0000;
      coeffs_in_data_log_force[5746] <= 16'h0000;
      coeffs_in_data_log_force[5747] <= 16'h0000;
      coeffs_in_data_log_force[5748] <= 16'h0000;
      coeffs_in_data_log_force[5749] <= 16'h0000;
      coeffs_in_data_log_force[5750] <= 16'h0000;
      coeffs_in_data_log_force[5751] <= 16'h0000;
      coeffs_in_data_log_force[5752] <= 16'h0000;
      coeffs_in_data_log_force[5753] <= 16'h0000;
      coeffs_in_data_log_force[5754] <= 16'h0000;
      coeffs_in_data_log_force[5755] <= 16'h0000;
      coeffs_in_data_log_force[5756] <= 16'h0000;
      coeffs_in_data_log_force[5757] <= 16'h0000;
      coeffs_in_data_log_force[5758] <= 16'h0000;
      coeffs_in_data_log_force[5759] <= 16'h0000;
      coeffs_in_data_log_force[5760] <= 16'h0000;
      coeffs_in_data_log_force[5761] <= 16'h0000;
      coeffs_in_data_log_force[5762] <= 16'h0000;
      coeffs_in_data_log_force[5763] <= 16'h0000;
      coeffs_in_data_log_force[5764] <= 16'h0000;
      coeffs_in_data_log_force[5765] <= 16'h0000;
      coeffs_in_data_log_force[5766] <= 16'h0000;
      coeffs_in_data_log_force[5767] <= 16'h0000;
      coeffs_in_data_log_force[5768] <= 16'h0000;
      coeffs_in_data_log_force[5769] <= 16'h0000;
      coeffs_in_data_log_force[5770] <= 16'h0000;
      coeffs_in_data_log_force[5771] <= 16'h0000;
      coeffs_in_data_log_force[5772] <= 16'h0000;
      coeffs_in_data_log_force[5773] <= 16'h0000;
      coeffs_in_data_log_force[5774] <= 16'h0000;
      coeffs_in_data_log_force[5775] <= 16'h0000;
      coeffs_in_data_log_force[5776] <= 16'h0000;
      coeffs_in_data_log_force[5777] <= 16'h0000;
      coeffs_in_data_log_force[5778] <= 16'h0000;
      coeffs_in_data_log_force[5779] <= 16'h0000;
      coeffs_in_data_log_force[5780] <= 16'h0000;
      coeffs_in_data_log_force[5781] <= 16'h0000;
      coeffs_in_data_log_force[5782] <= 16'h0000;
      coeffs_in_data_log_force[5783] <= 16'h0000;
      coeffs_in_data_log_force[5784] <= 16'h0000;
      coeffs_in_data_log_force[5785] <= 16'h0000;
      coeffs_in_data_log_force[5786] <= 16'h0000;
      coeffs_in_data_log_force[5787] <= 16'h0000;
      coeffs_in_data_log_force[5788] <= 16'h0000;
      coeffs_in_data_log_force[5789] <= 16'h0000;
      coeffs_in_data_log_force[5790] <= 16'h0000;
      coeffs_in_data_log_force[5791] <= 16'h0000;
      coeffs_in_data_log_force[5792] <= 16'h0000;
      coeffs_in_data_log_force[5793] <= 16'h0000;
      coeffs_in_data_log_force[5794] <= 16'h0000;
      coeffs_in_data_log_force[5795] <= 16'h0000;
      coeffs_in_data_log_force[5796] <= 16'h0000;
      coeffs_in_data_log_force[5797] <= 16'h0000;
      coeffs_in_data_log_force[5798] <= 16'h0000;
      coeffs_in_data_log_force[5799] <= 16'h0000;
      coeffs_in_data_log_force[5800] <= 16'h0000;
      coeffs_in_data_log_force[5801] <= 16'h0000;
      coeffs_in_data_log_force[5802] <= 16'h0000;
      coeffs_in_data_log_force[5803] <= 16'h0000;
      coeffs_in_data_log_force[5804] <= 16'h0000;
      coeffs_in_data_log_force[5805] <= 16'h0000;
      coeffs_in_data_log_force[5806] <= 16'h0000;
      coeffs_in_data_log_force[5807] <= 16'h0000;
      coeffs_in_data_log_force[5808] <= 16'h0000;
      coeffs_in_data_log_force[5809] <= 16'h0000;
      coeffs_in_data_log_force[5810] <= 16'h0000;
      coeffs_in_data_log_force[5811] <= 16'h0000;
      coeffs_in_data_log_force[5812] <= 16'h0000;
      coeffs_in_data_log_force[5813] <= 16'h0000;
      coeffs_in_data_log_force[5814] <= 16'h0000;
      coeffs_in_data_log_force[5815] <= 16'h0000;
      coeffs_in_data_log_force[5816] <= 16'h0000;
      coeffs_in_data_log_force[5817] <= 16'h0000;
      coeffs_in_data_log_force[5818] <= 16'h0000;
      coeffs_in_data_log_force[5819] <= 16'h0000;
      coeffs_in_data_log_force[5820] <= 16'h0000;
      coeffs_in_data_log_force[5821] <= 16'h0000;
      coeffs_in_data_log_force[5822] <= 16'h0000;
      coeffs_in_data_log_force[5823] <= 16'h0000;
      coeffs_in_data_log_force[5824] <= 16'h0000;
      coeffs_in_data_log_force[5825] <= 16'h0000;
      coeffs_in_data_log_force[5826] <= 16'h0000;
      coeffs_in_data_log_force[5827] <= 16'h0000;
      coeffs_in_data_log_force[5828] <= 16'h0000;
      coeffs_in_data_log_force[5829] <= 16'h0000;
      coeffs_in_data_log_force[5830] <= 16'h0000;
      coeffs_in_data_log_force[5831] <= 16'h0000;
      coeffs_in_data_log_force[5832] <= 16'h0000;
      coeffs_in_data_log_force[5833] <= 16'h0000;
      coeffs_in_data_log_force[5834] <= 16'h0000;
      coeffs_in_data_log_force[5835] <= 16'h0000;
      coeffs_in_data_log_force[5836] <= 16'h0000;
      coeffs_in_data_log_force[5837] <= 16'h0000;
      coeffs_in_data_log_force[5838] <= 16'h0000;
      coeffs_in_data_log_force[5839] <= 16'h0000;
      coeffs_in_data_log_force[5840] <= 16'h0000;
      coeffs_in_data_log_force[5841] <= 16'h0000;
      coeffs_in_data_log_force[5842] <= 16'h0000;
      coeffs_in_data_log_force[5843] <= 16'h0000;
      coeffs_in_data_log_force[5844] <= 16'h0000;
      coeffs_in_data_log_force[5845] <= 16'h0000;
      coeffs_in_data_log_force[5846] <= 16'h0000;
      coeffs_in_data_log_force[5847] <= 16'h0000;
      coeffs_in_data_log_force[5848] <= 16'h0000;
      coeffs_in_data_log_force[5849] <= 16'h0000;
      coeffs_in_data_log_force[5850] <= 16'h0000;
      coeffs_in_data_log_force[5851] <= 16'h0000;
      coeffs_in_data_log_force[5852] <= 16'h0000;
      coeffs_in_data_log_force[5853] <= 16'h0000;
      coeffs_in_data_log_force[5854] <= 16'h0000;
      coeffs_in_data_log_force[5855] <= 16'h0000;
      coeffs_in_data_log_force[5856] <= 16'h0000;
      coeffs_in_data_log_force[5857] <= 16'h0000;
      coeffs_in_data_log_force[5858] <= 16'h0000;
      coeffs_in_data_log_force[5859] <= 16'h0000;
      coeffs_in_data_log_force[5860] <= 16'h0000;
      coeffs_in_data_log_force[5861] <= 16'h0000;
      coeffs_in_data_log_force[5862] <= 16'h0000;
      coeffs_in_data_log_force[5863] <= 16'h0000;
      coeffs_in_data_log_force[5864] <= 16'h0000;
      coeffs_in_data_log_force[5865] <= 16'h0000;
      coeffs_in_data_log_force[5866] <= 16'h0000;
      coeffs_in_data_log_force[5867] <= 16'h0000;
      coeffs_in_data_log_force[5868] <= 16'h0000;
      coeffs_in_data_log_force[5869] <= 16'h0000;
      coeffs_in_data_log_force[5870] <= 16'h0000;
      coeffs_in_data_log_force[5871] <= 16'h0000;
      coeffs_in_data_log_force[5872] <= 16'h0000;
      coeffs_in_data_log_force[5873] <= 16'h0000;
      coeffs_in_data_log_force[5874] <= 16'h0000;
      coeffs_in_data_log_force[5875] <= 16'h0000;
      coeffs_in_data_log_force[5876] <= 16'h0000;
      coeffs_in_data_log_force[5877] <= 16'h0000;
      coeffs_in_data_log_force[5878] <= 16'h0000;
      coeffs_in_data_log_force[5879] <= 16'h0000;
      coeffs_in_data_log_force[5880] <= 16'h0000;
      coeffs_in_data_log_force[5881] <= 16'h0000;
      coeffs_in_data_log_force[5882] <= 16'h0000;
      coeffs_in_data_log_force[5883] <= 16'h0000;
      coeffs_in_data_log_force[5884] <= 16'h0000;
      coeffs_in_data_log_force[5885] <= 16'h0000;
      coeffs_in_data_log_force[5886] <= 16'h0000;
      coeffs_in_data_log_force[5887] <= 16'h0000;
      coeffs_in_data_log_force[5888] <= 16'h0000;
      coeffs_in_data_log_force[5889] <= 16'h0000;
      coeffs_in_data_log_force[5890] <= 16'h0000;
      coeffs_in_data_log_force[5891] <= 16'h0000;
      coeffs_in_data_log_force[5892] <= 16'h0000;
      coeffs_in_data_log_force[5893] <= 16'h0000;
      coeffs_in_data_log_force[5894] <= 16'h0000;
      coeffs_in_data_log_force[5895] <= 16'h0000;
      coeffs_in_data_log_force[5896] <= 16'h0000;
      coeffs_in_data_log_force[5897] <= 16'h0000;
      coeffs_in_data_log_force[5898] <= 16'h0000;
      coeffs_in_data_log_force[5899] <= 16'h0000;
      coeffs_in_data_log_force[5900] <= 16'h0000;
      coeffs_in_data_log_force[5901] <= 16'h0000;
      coeffs_in_data_log_force[5902] <= 16'h0000;
      coeffs_in_data_log_force[5903] <= 16'h0000;
      coeffs_in_data_log_force[5904] <= 16'h0000;
      coeffs_in_data_log_force[5905] <= 16'h0000;
      coeffs_in_data_log_force[5906] <= 16'h0000;
      coeffs_in_data_log_force[5907] <= 16'h0000;
      coeffs_in_data_log_force[5908] <= 16'h0000;
      coeffs_in_data_log_force[5909] <= 16'h0000;
      coeffs_in_data_log_force[5910] <= 16'h0000;
      coeffs_in_data_log_force[5911] <= 16'h0000;
      coeffs_in_data_log_force[5912] <= 16'h0000;
      coeffs_in_data_log_force[5913] <= 16'h0000;
      coeffs_in_data_log_force[5914] <= 16'h0000;
      coeffs_in_data_log_force[5915] <= 16'h0000;
      coeffs_in_data_log_force[5916] <= 16'h0000;
      coeffs_in_data_log_force[5917] <= 16'h0000;
      coeffs_in_data_log_force[5918] <= 16'h0000;
      coeffs_in_data_log_force[5919] <= 16'h0000;
      coeffs_in_data_log_force[5920] <= 16'h0000;
      coeffs_in_data_log_force[5921] <= 16'h0000;
      coeffs_in_data_log_force[5922] <= 16'h0000;
      coeffs_in_data_log_force[5923] <= 16'h0000;
      coeffs_in_data_log_force[5924] <= 16'h0000;
      coeffs_in_data_log_force[5925] <= 16'h0000;
      coeffs_in_data_log_force[5926] <= 16'h0000;
      coeffs_in_data_log_force[5927] <= 16'h0000;
      coeffs_in_data_log_force[5928] <= 16'h0000;
      coeffs_in_data_log_force[5929] <= 16'h0000;
      coeffs_in_data_log_force[5930] <= 16'h0000;
      coeffs_in_data_log_force[5931] <= 16'h0000;
      coeffs_in_data_log_force[5932] <= 16'h0000;
      coeffs_in_data_log_force[5933] <= 16'h0000;
      coeffs_in_data_log_force[5934] <= 16'h0000;
      coeffs_in_data_log_force[5935] <= 16'h0000;
      coeffs_in_data_log_force[5936] <= 16'h0000;
      coeffs_in_data_log_force[5937] <= 16'h0000;
      coeffs_in_data_log_force[5938] <= 16'h0000;
      coeffs_in_data_log_force[5939] <= 16'h0000;
      coeffs_in_data_log_force[5940] <= 16'h0000;
      coeffs_in_data_log_force[5941] <= 16'h0000;
      coeffs_in_data_log_force[5942] <= 16'h0000;
      coeffs_in_data_log_force[5943] <= 16'h0000;
      coeffs_in_data_log_force[5944] <= 16'h0000;
      coeffs_in_data_log_force[5945] <= 16'h0000;
      coeffs_in_data_log_force[5946] <= 16'h0000;
      coeffs_in_data_log_force[5947] <= 16'h0000;
      coeffs_in_data_log_force[5948] <= 16'h0000;
      coeffs_in_data_log_force[5949] <= 16'h0000;
      coeffs_in_data_log_force[5950] <= 16'h0000;
      coeffs_in_data_log_force[5951] <= 16'h0000;
      coeffs_in_data_log_force[5952] <= 16'h0000;
      coeffs_in_data_log_force[5953] <= 16'h0000;
      coeffs_in_data_log_force[5954] <= 16'h0000;
      coeffs_in_data_log_force[5955] <= 16'h0000;
      coeffs_in_data_log_force[5956] <= 16'h0000;
      coeffs_in_data_log_force[5957] <= 16'h0000;
      coeffs_in_data_log_force[5958] <= 16'h0000;
      coeffs_in_data_log_force[5959] <= 16'h0000;
      coeffs_in_data_log_force[5960] <= 16'h0000;
      coeffs_in_data_log_force[5961] <= 16'h0000;
      coeffs_in_data_log_force[5962] <= 16'h0000;
      coeffs_in_data_log_force[5963] <= 16'h0000;
      coeffs_in_data_log_force[5964] <= 16'h0000;
      coeffs_in_data_log_force[5965] <= 16'h0000;
      coeffs_in_data_log_force[5966] <= 16'h0000;
      coeffs_in_data_log_force[5967] <= 16'h0000;
      coeffs_in_data_log_force[5968] <= 16'h0000;
      coeffs_in_data_log_force[5969] <= 16'h0000;
      coeffs_in_data_log_force[5970] <= 16'h0000;
      coeffs_in_data_log_force[5971] <= 16'h0000;
      coeffs_in_data_log_force[5972] <= 16'h0000;
      coeffs_in_data_log_force[5973] <= 16'h0000;
      coeffs_in_data_log_force[5974] <= 16'h0000;
      coeffs_in_data_log_force[5975] <= 16'h0000;
      coeffs_in_data_log_force[5976] <= 16'h0000;
      coeffs_in_data_log_force[5977] <= 16'h0000;
      coeffs_in_data_log_force[5978] <= 16'h0000;
      coeffs_in_data_log_force[5979] <= 16'h0000;
      coeffs_in_data_log_force[5980] <= 16'h0000;
      coeffs_in_data_log_force[5981] <= 16'h0000;
      coeffs_in_data_log_force[5982] <= 16'h0000;
      coeffs_in_data_log_force[5983] <= 16'h0000;
      coeffs_in_data_log_force[5984] <= 16'h0000;
      coeffs_in_data_log_force[5985] <= 16'h0000;
      coeffs_in_data_log_force[5986] <= 16'h0000;
      coeffs_in_data_log_force[5987] <= 16'h0000;
      coeffs_in_data_log_force[5988] <= 16'h0000;
      coeffs_in_data_log_force[5989] <= 16'h0000;
      coeffs_in_data_log_force[5990] <= 16'h0000;
      coeffs_in_data_log_force[5991] <= 16'h0000;
      coeffs_in_data_log_force[5992] <= 16'h0000;
      coeffs_in_data_log_force[5993] <= 16'h0000;
      coeffs_in_data_log_force[5994] <= 16'h0000;
      coeffs_in_data_log_force[5995] <= 16'h0000;
      coeffs_in_data_log_force[5996] <= 16'h0000;
      coeffs_in_data_log_force[5997] <= 16'h0000;
      coeffs_in_data_log_force[5998] <= 16'h0000;
      coeffs_in_data_log_force[5999] <= 16'h0000;
      coeffs_in_data_log_force[6000] <= 16'h0000;
      coeffs_in_data_log_force[6001] <= 16'h0000;
      coeffs_in_data_log_force[6002] <= 16'h0000;
      coeffs_in_data_log_force[6003] <= 16'h0000;
      coeffs_in_data_log_force[6004] <= 16'h0000;
      coeffs_in_data_log_force[6005] <= 16'h0000;
      coeffs_in_data_log_force[6006] <= 16'h0000;
      coeffs_in_data_log_force[6007] <= 16'h0000;
      coeffs_in_data_log_force[6008] <= 16'h0000;
      coeffs_in_data_log_force[6009] <= 16'h0000;
      coeffs_in_data_log_force[6010] <= 16'h0000;
      coeffs_in_data_log_force[6011] <= 16'h0000;
      coeffs_in_data_log_force[6012] <= 16'h0000;
      coeffs_in_data_log_force[6013] <= 16'h0000;
      coeffs_in_data_log_force[6014] <= 16'h0000;
      coeffs_in_data_log_force[6015] <= 16'h0000;
      coeffs_in_data_log_force[6016] <= 16'h0000;
      coeffs_in_data_log_force[6017] <= 16'h0000;
      coeffs_in_data_log_force[6018] <= 16'h0000;
      coeffs_in_data_log_force[6019] <= 16'h0000;
      coeffs_in_data_log_force[6020] <= 16'h0000;
      coeffs_in_data_log_force[6021] <= 16'h0000;
      coeffs_in_data_log_force[6022] <= 16'h0000;
      coeffs_in_data_log_force[6023] <= 16'h0000;
      coeffs_in_data_log_force[6024] <= 16'h0000;
      coeffs_in_data_log_force[6025] <= 16'h0000;
      coeffs_in_data_log_force[6026] <= 16'h0000;
      coeffs_in_data_log_force[6027] <= 16'h0000;
      coeffs_in_data_log_force[6028] <= 16'h0000;
      coeffs_in_data_log_force[6029] <= 16'h0000;
      coeffs_in_data_log_force[6030] <= 16'h0000;
      coeffs_in_data_log_force[6031] <= 16'h0000;
      coeffs_in_data_log_force[6032] <= 16'h0000;
      coeffs_in_data_log_force[6033] <= 16'h0000;
      coeffs_in_data_log_force[6034] <= 16'h0000;
      coeffs_in_data_log_force[6035] <= 16'h0000;
      coeffs_in_data_log_force[6036] <= 16'h0000;
      coeffs_in_data_log_force[6037] <= 16'h0000;
      coeffs_in_data_log_force[6038] <= 16'h0000;
      coeffs_in_data_log_force[6039] <= 16'h0000;
      coeffs_in_data_log_force[6040] <= 16'h0000;
      coeffs_in_data_log_force[6041] <= 16'h0000;
      coeffs_in_data_log_force[6042] <= 16'h0000;
      coeffs_in_data_log_force[6043] <= 16'h0000;
      coeffs_in_data_log_force[6044] <= 16'h0000;
      coeffs_in_data_log_force[6045] <= 16'h0000;
      coeffs_in_data_log_force[6046] <= 16'h0000;
      coeffs_in_data_log_force[6047] <= 16'h0000;
      coeffs_in_data_log_force[6048] <= 16'h0000;
      coeffs_in_data_log_force[6049] <= 16'h0000;
      coeffs_in_data_log_force[6050] <= 16'h0000;
      coeffs_in_data_log_force[6051] <= 16'h0000;
      coeffs_in_data_log_force[6052] <= 16'h0000;
      coeffs_in_data_log_force[6053] <= 16'h0000;
      coeffs_in_data_log_force[6054] <= 16'h0000;
      coeffs_in_data_log_force[6055] <= 16'h0000;
      coeffs_in_data_log_force[6056] <= 16'h0000;
      coeffs_in_data_log_force[6057] <= 16'h0000;
      coeffs_in_data_log_force[6058] <= 16'h0000;
      coeffs_in_data_log_force[6059] <= 16'h0000;
      coeffs_in_data_log_force[6060] <= 16'h0000;
      coeffs_in_data_log_force[6061] <= 16'h0000;
      coeffs_in_data_log_force[6062] <= 16'h0000;
      coeffs_in_data_log_force[6063] <= 16'h0000;
      coeffs_in_data_log_force[6064] <= 16'h0000;
      coeffs_in_data_log_force[6065] <= 16'h0000;
      coeffs_in_data_log_force[6066] <= 16'h0000;
      coeffs_in_data_log_force[6067] <= 16'h0000;
      coeffs_in_data_log_force[6068] <= 16'h0000;
      coeffs_in_data_log_force[6069] <= 16'h0000;
      coeffs_in_data_log_force[6070] <= 16'h0000;
      coeffs_in_data_log_force[6071] <= 16'h0000;
      coeffs_in_data_log_force[6072] <= 16'h0000;
      coeffs_in_data_log_force[6073] <= 16'h0000;
      coeffs_in_data_log_force[6074] <= 16'h0000;
      coeffs_in_data_log_force[6075] <= 16'h0000;
      coeffs_in_data_log_force[6076] <= 16'h0000;
      coeffs_in_data_log_force[6077] <= 16'h0000;
      coeffs_in_data_log_force[6078] <= 16'h0000;
      coeffs_in_data_log_force[6079] <= 16'h0000;
      coeffs_in_data_log_force[6080] <= 16'h0000;
      coeffs_in_data_log_force[6081] <= 16'h0000;
      coeffs_in_data_log_force[6082] <= 16'h0000;
      coeffs_in_data_log_force[6083] <= 16'h0000;
      coeffs_in_data_log_force[6084] <= 16'h0000;
      coeffs_in_data_log_force[6085] <= 16'h0000;
      coeffs_in_data_log_force[6086] <= 16'h0000;
      coeffs_in_data_log_force[6087] <= 16'h0000;
      coeffs_in_data_log_force[6088] <= 16'h0000;
      coeffs_in_data_log_force[6089] <= 16'h0000;
      coeffs_in_data_log_force[6090] <= 16'h0000;
      coeffs_in_data_log_force[6091] <= 16'h0000;
      coeffs_in_data_log_force[6092] <= 16'h0000;
      coeffs_in_data_log_force[6093] <= 16'h0000;
      coeffs_in_data_log_force[6094] <= 16'h0000;
      coeffs_in_data_log_force[6095] <= 16'h0000;
      coeffs_in_data_log_force[6096] <= 16'h0000;
      coeffs_in_data_log_force[6097] <= 16'h0000;
      coeffs_in_data_log_force[6098] <= 16'h0000;
      coeffs_in_data_log_force[6099] <= 16'h0000;
      coeffs_in_data_log_force[6100] <= 16'h0000;
      coeffs_in_data_log_force[6101] <= 16'h0000;
      coeffs_in_data_log_force[6102] <= 16'h0000;
      coeffs_in_data_log_force[6103] <= 16'h0000;
      coeffs_in_data_log_force[6104] <= 16'h0000;
      coeffs_in_data_log_force[6105] <= 16'h0000;
      coeffs_in_data_log_force[6106] <= 16'h0000;
      coeffs_in_data_log_force[6107] <= 16'h0000;
      coeffs_in_data_log_force[6108] <= 16'h0000;
      coeffs_in_data_log_force[6109] <= 16'h0000;
      coeffs_in_data_log_force[6110] <= 16'h0000;
      coeffs_in_data_log_force[6111] <= 16'h0000;
      coeffs_in_data_log_force[6112] <= 16'h0000;
      coeffs_in_data_log_force[6113] <= 16'h0000;
      coeffs_in_data_log_force[6114] <= 16'h0000;
      coeffs_in_data_log_force[6115] <= 16'h0000;
      coeffs_in_data_log_force[6116] <= 16'h0000;
      coeffs_in_data_log_force[6117] <= 16'h0000;
      coeffs_in_data_log_force[6118] <= 16'h0000;
      coeffs_in_data_log_force[6119] <= 16'h0000;
      coeffs_in_data_log_force[6120] <= 16'h0000;
      coeffs_in_data_log_force[6121] <= 16'h0000;
      coeffs_in_data_log_force[6122] <= 16'h0000;
      coeffs_in_data_log_force[6123] <= 16'h0000;
      coeffs_in_data_log_force[6124] <= 16'h0000;
      coeffs_in_data_log_force[6125] <= 16'h0000;
      coeffs_in_data_log_force[6126] <= 16'h0000;
      coeffs_in_data_log_force[6127] <= 16'h0000;
      coeffs_in_data_log_force[6128] <= 16'h0000;
      coeffs_in_data_log_force[6129] <= 16'h0000;
      coeffs_in_data_log_force[6130] <= 16'h0000;
      coeffs_in_data_log_force[6131] <= 16'h0000;
      coeffs_in_data_log_force[6132] <= 16'h0000;
      coeffs_in_data_log_force[6133] <= 16'h0000;
      coeffs_in_data_log_force[6134] <= 16'h0000;
      coeffs_in_data_log_force[6135] <= 16'h0000;
      coeffs_in_data_log_force[6136] <= 16'h0000;
      coeffs_in_data_log_force[6137] <= 16'h0000;
      coeffs_in_data_log_force[6138] <= 16'h0000;
      coeffs_in_data_log_force[6139] <= 16'h0000;
      coeffs_in_data_log_force[6140] <= 16'h0000;
      coeffs_in_data_log_force[6141] <= 16'h0000;
      coeffs_in_data_log_force[6142] <= 16'h0000;
      coeffs_in_data_log_force[6143] <= 16'h0000;
      coeffs_in_data_log_force[6144] <= 16'h0000;
      coeffs_in_data_log_force[6145] <= 16'h0000;
      coeffs_in_data_log_force[6146] <= 16'h0000;
      coeffs_in_data_log_force[6147] <= 16'h0000;
      coeffs_in_data_log_force[6148] <= 16'h0000;
      coeffs_in_data_log_force[6149] <= 16'h0000;
      coeffs_in_data_log_force[6150] <= 16'h0000;
      coeffs_in_data_log_force[6151] <= 16'h0000;
      coeffs_in_data_log_force[6152] <= 16'h0000;
      coeffs_in_data_log_force[6153] <= 16'h0000;
      coeffs_in_data_log_force[6154] <= 16'h0000;
      coeffs_in_data_log_force[6155] <= 16'h0000;
      coeffs_in_data_log_force[6156] <= 16'h0000;
      coeffs_in_data_log_force[6157] <= 16'h0000;
      coeffs_in_data_log_force[6158] <= 16'h0000;
      coeffs_in_data_log_force[6159] <= 16'h0000;
      coeffs_in_data_log_force[6160] <= 16'h0000;
      coeffs_in_data_log_force[6161] <= 16'h0000;
      coeffs_in_data_log_force[6162] <= 16'h0000;
      coeffs_in_data_log_force[6163] <= 16'h0000;
      coeffs_in_data_log_force[6164] <= 16'h0000;
      coeffs_in_data_log_force[6165] <= 16'h0000;
      coeffs_in_data_log_force[6166] <= 16'h0000;
      coeffs_in_data_log_force[6167] <= 16'h0000;
      coeffs_in_data_log_force[6168] <= 16'h0000;
      coeffs_in_data_log_force[6169] <= 16'h0000;
      coeffs_in_data_log_force[6170] <= 16'h0000;
      coeffs_in_data_log_force[6171] <= 16'h0000;
      coeffs_in_data_log_force[6172] <= 16'h0000;
      coeffs_in_data_log_force[6173] <= 16'h0000;
      coeffs_in_data_log_force[6174] <= 16'h0000;
      coeffs_in_data_log_force[6175] <= 16'h0000;
      coeffs_in_data_log_force[6176] <= 16'h0000;
      coeffs_in_data_log_force[6177] <= 16'h0000;
      coeffs_in_data_log_force[6178] <= 16'h0000;
      coeffs_in_data_log_force[6179] <= 16'h0000;
      coeffs_in_data_log_force[6180] <= 16'h0000;
      coeffs_in_data_log_force[6181] <= 16'h0000;
      coeffs_in_data_log_force[6182] <= 16'h0000;
      coeffs_in_data_log_force[6183] <= 16'h0000;
      coeffs_in_data_log_force[6184] <= 16'h0000;
      coeffs_in_data_log_force[6185] <= 16'h0000;
      coeffs_in_data_log_force[6186] <= 16'h0000;
      coeffs_in_data_log_force[6187] <= 16'h0000;
      coeffs_in_data_log_force[6188] <= 16'h0000;
      coeffs_in_data_log_force[6189] <= 16'h0000;
      coeffs_in_data_log_force[6190] <= 16'h0000;
      coeffs_in_data_log_force[6191] <= 16'h0000;
      coeffs_in_data_log_force[6192] <= 16'h0000;
      coeffs_in_data_log_force[6193] <= 16'h0000;
      coeffs_in_data_log_force[6194] <= 16'h0000;
      coeffs_in_data_log_force[6195] <= 16'h0000;
      coeffs_in_data_log_force[6196] <= 16'h0000;
      coeffs_in_data_log_force[6197] <= 16'h0000;
      coeffs_in_data_log_force[6198] <= 16'h0000;
      coeffs_in_data_log_force[6199] <= 16'h0000;
      coeffs_in_data_log_force[6200] <= 16'h0000;
      coeffs_in_data_log_force[6201] <= 16'h0000;
      coeffs_in_data_log_force[6202] <= 16'h0000;
      coeffs_in_data_log_force[6203] <= 16'h0000;
      coeffs_in_data_log_force[6204] <= 16'h0000;
      coeffs_in_data_log_force[6205] <= 16'h0000;
      coeffs_in_data_log_force[6206] <= 16'h0000;
      coeffs_in_data_log_force[6207] <= 16'h0000;
      coeffs_in_data_log_force[6208] <= 16'h0000;
      coeffs_in_data_log_force[6209] <= 16'h0000;
      coeffs_in_data_log_force[6210] <= 16'h0000;
      coeffs_in_data_log_force[6211] <= 16'h0000;
      coeffs_in_data_log_force[6212] <= 16'h0000;
      coeffs_in_data_log_force[6213] <= 16'h0000;
      coeffs_in_data_log_force[6214] <= 16'h0000;
      coeffs_in_data_log_force[6215] <= 16'h0000;
      coeffs_in_data_log_force[6216] <= 16'h0000;
      coeffs_in_data_log_force[6217] <= 16'h0000;
      coeffs_in_data_log_force[6218] <= 16'h0000;
      coeffs_in_data_log_force[6219] <= 16'h0000;
      coeffs_in_data_log_force[6220] <= 16'h0000;
      coeffs_in_data_log_force[6221] <= 16'h0000;
      coeffs_in_data_log_force[6222] <= 16'h0000;
      coeffs_in_data_log_force[6223] <= 16'h0000;
      coeffs_in_data_log_force[6224] <= 16'h0000;
      coeffs_in_data_log_force[6225] <= 16'h0000;
      coeffs_in_data_log_force[6226] <= 16'h0000;
      coeffs_in_data_log_force[6227] <= 16'h0000;
      coeffs_in_data_log_force[6228] <= 16'h0000;
      coeffs_in_data_log_force[6229] <= 16'h0000;
      coeffs_in_data_log_force[6230] <= 16'h0000;
      coeffs_in_data_log_force[6231] <= 16'h0000;
      coeffs_in_data_log_force[6232] <= 16'h0000;
      coeffs_in_data_log_force[6233] <= 16'h0000;
      coeffs_in_data_log_force[6234] <= 16'h0000;
      coeffs_in_data_log_force[6235] <= 16'h0000;
      coeffs_in_data_log_force[6236] <= 16'h0000;
      coeffs_in_data_log_force[6237] <= 16'h0000;
      coeffs_in_data_log_force[6238] <= 16'h0000;
      coeffs_in_data_log_force[6239] <= 16'h0000;
      coeffs_in_data_log_force[6240] <= 16'h0000;
      coeffs_in_data_log_force[6241] <= 16'h0000;
      coeffs_in_data_log_force[6242] <= 16'h0000;
      coeffs_in_data_log_force[6243] <= 16'h0000;
      coeffs_in_data_log_force[6244] <= 16'h0000;
      coeffs_in_data_log_force[6245] <= 16'h0000;
      coeffs_in_data_log_force[6246] <= 16'h0000;
      coeffs_in_data_log_force[6247] <= 16'h0000;
      coeffs_in_data_log_force[6248] <= 16'h0000;
      coeffs_in_data_log_force[6249] <= 16'h0000;
      coeffs_in_data_log_force[6250] <= 16'h0000;
      coeffs_in_data_log_force[6251] <= 16'h0000;
      coeffs_in_data_log_force[6252] <= 16'h0000;
      coeffs_in_data_log_force[6253] <= 16'h0000;
      coeffs_in_data_log_force[6254] <= 16'h0000;
      coeffs_in_data_log_force[6255] <= 16'h0000;
      coeffs_in_data_log_force[6256] <= 16'h0000;
      coeffs_in_data_log_force[6257] <= 16'h0000;
      coeffs_in_data_log_force[6258] <= 16'h0000;
      coeffs_in_data_log_force[6259] <= 16'h0000;
      coeffs_in_data_log_force[6260] <= 16'h0000;
      coeffs_in_data_log_force[6261] <= 16'h0000;
      coeffs_in_data_log_force[6262] <= 16'h0000;
      coeffs_in_data_log_force[6263] <= 16'h0000;
      coeffs_in_data_log_force[6264] <= 16'h0000;
      coeffs_in_data_log_force[6265] <= 16'h0000;
      coeffs_in_data_log_force[6266] <= 16'h0000;
      coeffs_in_data_log_force[6267] <= 16'h0000;
      coeffs_in_data_log_force[6268] <= 16'h0000;
      coeffs_in_data_log_force[6269] <= 16'h0000;
      coeffs_in_data_log_force[6270] <= 16'h0000;
      coeffs_in_data_log_force[6271] <= 16'h0000;
      coeffs_in_data_log_force[6272] <= 16'h0000;
      coeffs_in_data_log_force[6273] <= 16'h0000;
      coeffs_in_data_log_force[6274] <= 16'h0000;
      coeffs_in_data_log_force[6275] <= 16'h0000;
      coeffs_in_data_log_force[6276] <= 16'h0000;
      coeffs_in_data_log_force[6277] <= 16'h0000;
      coeffs_in_data_log_force[6278] <= 16'h0000;
      coeffs_in_data_log_force[6279] <= 16'h0000;
      coeffs_in_data_log_force[6280] <= 16'h0000;
      coeffs_in_data_log_force[6281] <= 16'h0000;
      coeffs_in_data_log_force[6282] <= 16'h0000;
      coeffs_in_data_log_force[6283] <= 16'h0000;
      coeffs_in_data_log_force[6284] <= 16'h0000;
      coeffs_in_data_log_force[6285] <= 16'h0000;
      coeffs_in_data_log_force[6286] <= 16'h0000;
      coeffs_in_data_log_force[6287] <= 16'h0000;
      coeffs_in_data_log_force[6288] <= 16'h0000;
      coeffs_in_data_log_force[6289] <= 16'h0000;
      coeffs_in_data_log_force[6290] <= 16'h0000;
      coeffs_in_data_log_force[6291] <= 16'h0000;
      coeffs_in_data_log_force[6292] <= 16'h0000;
      coeffs_in_data_log_force[6293] <= 16'h0000;
      coeffs_in_data_log_force[6294] <= 16'h0000;
      coeffs_in_data_log_force[6295] <= 16'h0000;
      coeffs_in_data_log_force[6296] <= 16'h0000;
      coeffs_in_data_log_force[6297] <= 16'h0000;
      coeffs_in_data_log_force[6298] <= 16'h0000;
      coeffs_in_data_log_force[6299] <= 16'h0000;
      coeffs_in_data_log_force[6300] <= 16'h0000;
      coeffs_in_data_log_force[6301] <= 16'h0000;
      coeffs_in_data_log_force[6302] <= 16'h0000;
      coeffs_in_data_log_force[6303] <= 16'h0000;
      coeffs_in_data_log_force[6304] <= 16'h0000;
      coeffs_in_data_log_force[6305] <= 16'h0000;
      coeffs_in_data_log_force[6306] <= 16'h0000;
      coeffs_in_data_log_force[6307] <= 16'h0000;
      coeffs_in_data_log_force[6308] <= 16'h0000;
      coeffs_in_data_log_force[6309] <= 16'h0000;
      coeffs_in_data_log_force[6310] <= 16'h0000;
      coeffs_in_data_log_force[6311] <= 16'h0000;
      coeffs_in_data_log_force[6312] <= 16'h0000;
      coeffs_in_data_log_force[6313] <= 16'h0000;
      coeffs_in_data_log_force[6314] <= 16'h0000;
      coeffs_in_data_log_force[6315] <= 16'h0000;
      coeffs_in_data_log_force[6316] <= 16'h0000;
      coeffs_in_data_log_force[6317] <= 16'h0000;
      coeffs_in_data_log_force[6318] <= 16'h0000;
      coeffs_in_data_log_force[6319] <= 16'h0000;
      coeffs_in_data_log_force[6320] <= 16'h0000;
      coeffs_in_data_log_force[6321] <= 16'h0000;
      coeffs_in_data_log_force[6322] <= 16'h0000;
      coeffs_in_data_log_force[6323] <= 16'h0000;
      coeffs_in_data_log_force[6324] <= 16'h0000;
      coeffs_in_data_log_force[6325] <= 16'h0000;
      coeffs_in_data_log_force[6326] <= 16'h0000;
      coeffs_in_data_log_force[6327] <= 16'h0000;
      coeffs_in_data_log_force[6328] <= 16'h0000;
      coeffs_in_data_log_force[6329] <= 16'h0000;
      coeffs_in_data_log_force[6330] <= 16'h0000;
      coeffs_in_data_log_force[6331] <= 16'h0000;
      coeffs_in_data_log_force[6332] <= 16'h0000;
      coeffs_in_data_log_force[6333] <= 16'h0000;
      coeffs_in_data_log_force[6334] <= 16'h0000;
      coeffs_in_data_log_force[6335] <= 16'h0000;
      coeffs_in_data_log_force[6336] <= 16'h0000;
      coeffs_in_data_log_force[6337] <= 16'h0000;
      coeffs_in_data_log_force[6338] <= 16'h0000;
      coeffs_in_data_log_force[6339] <= 16'h0000;
      coeffs_in_data_log_force[6340] <= 16'h0000;
      coeffs_in_data_log_force[6341] <= 16'h0000;
      coeffs_in_data_log_force[6342] <= 16'h0000;
      coeffs_in_data_log_force[6343] <= 16'h0000;
      coeffs_in_data_log_force[6344] <= 16'h0000;
      coeffs_in_data_log_force[6345] <= 16'h0000;
      coeffs_in_data_log_force[6346] <= 16'h0000;
      coeffs_in_data_log_force[6347] <= 16'h0000;
      coeffs_in_data_log_force[6348] <= 16'h0000;
      coeffs_in_data_log_force[6349] <= 16'h0000;
      coeffs_in_data_log_force[6350] <= 16'h0000;
      coeffs_in_data_log_force[6351] <= 16'h0000;
      coeffs_in_data_log_force[6352] <= 16'h0000;
      coeffs_in_data_log_force[6353] <= 16'h0000;
      coeffs_in_data_log_force[6354] <= 16'h0000;
      coeffs_in_data_log_force[6355] <= 16'h0000;
      coeffs_in_data_log_force[6356] <= 16'h0000;
      coeffs_in_data_log_force[6357] <= 16'h0000;
      coeffs_in_data_log_force[6358] <= 16'h0000;
      coeffs_in_data_log_force[6359] <= 16'h0000;
      coeffs_in_data_log_force[6360] <= 16'h0000;
      coeffs_in_data_log_force[6361] <= 16'h0000;
      coeffs_in_data_log_force[6362] <= 16'h0000;
      coeffs_in_data_log_force[6363] <= 16'h0000;
      coeffs_in_data_log_force[6364] <= 16'h0000;
      coeffs_in_data_log_force[6365] <= 16'h0000;
      coeffs_in_data_log_force[6366] <= 16'h0000;
      coeffs_in_data_log_force[6367] <= 16'h0000;
      coeffs_in_data_log_force[6368] <= 16'h0000;
      coeffs_in_data_log_force[6369] <= 16'h0000;
      coeffs_in_data_log_force[6370] <= 16'h0000;
      coeffs_in_data_log_force[6371] <= 16'h0000;
      coeffs_in_data_log_force[6372] <= 16'h0000;
      coeffs_in_data_log_force[6373] <= 16'h0000;
      coeffs_in_data_log_force[6374] <= 16'h0000;
      coeffs_in_data_log_force[6375] <= 16'h0000;
      coeffs_in_data_log_force[6376] <= 16'h0000;
      coeffs_in_data_log_force[6377] <= 16'h0000;
      coeffs_in_data_log_force[6378] <= 16'h0000;
      coeffs_in_data_log_force[6379] <= 16'h0000;
      coeffs_in_data_log_force[6380] <= 16'h0000;
      coeffs_in_data_log_force[6381] <= 16'h0000;
      coeffs_in_data_log_force[6382] <= 16'h0000;
      coeffs_in_data_log_force[6383] <= 16'h0000;
      coeffs_in_data_log_force[6384] <= 16'h0000;
      coeffs_in_data_log_force[6385] <= 16'h0000;
      coeffs_in_data_log_force[6386] <= 16'h0000;
      coeffs_in_data_log_force[6387] <= 16'h0000;
      coeffs_in_data_log_force[6388] <= 16'h0000;
      coeffs_in_data_log_force[6389] <= 16'h0000;
      coeffs_in_data_log_force[6390] <= 16'h0000;
      coeffs_in_data_log_force[6391] <= 16'h0000;
      coeffs_in_data_log_force[6392] <= 16'h0000;
      coeffs_in_data_log_force[6393] <= 16'h0000;
      coeffs_in_data_log_force[6394] <= 16'h0000;
      coeffs_in_data_log_force[6395] <= 16'h0000;
      coeffs_in_data_log_force[6396] <= 16'h0000;
      coeffs_in_data_log_force[6397] <= 16'h0000;
      coeffs_in_data_log_force[6398] <= 16'h0000;
      coeffs_in_data_log_force[6399] <= 16'h0000;
      coeffs_in_data_log_force[6400] <= 16'h0000;
      coeffs_in_data_log_force[6401] <= 16'h0000;
      coeffs_in_data_log_force[6402] <= 16'h0000;
      coeffs_in_data_log_force[6403] <= 16'h0000;
      coeffs_in_data_log_force[6404] <= 16'h0000;
      coeffs_in_data_log_force[6405] <= 16'h0000;
      coeffs_in_data_log_force[6406] <= 16'h0000;
      coeffs_in_data_log_force[6407] <= 16'h0000;
      coeffs_in_data_log_force[6408] <= 16'h0000;
      coeffs_in_data_log_force[6409] <= 16'h0000;
      coeffs_in_data_log_force[6410] <= 16'h0000;
      coeffs_in_data_log_force[6411] <= 16'h0000;
      coeffs_in_data_log_force[6412] <= 16'h0000;
      coeffs_in_data_log_force[6413] <= 16'h0000;
      coeffs_in_data_log_force[6414] <= 16'h0000;
      coeffs_in_data_log_force[6415] <= 16'h0000;
      coeffs_in_data_log_force[6416] <= 16'h0000;
      coeffs_in_data_log_force[6417] <= 16'h0000;
      coeffs_in_data_log_force[6418] <= 16'h0000;
      coeffs_in_data_log_force[6419] <= 16'h0000;
      coeffs_in_data_log_force[6420] <= 16'h0000;
      coeffs_in_data_log_force[6421] <= 16'h0000;
      coeffs_in_data_log_force[6422] <= 16'h0000;
      coeffs_in_data_log_force[6423] <= 16'h0000;
      coeffs_in_data_log_force[6424] <= 16'h0000;
      coeffs_in_data_log_force[6425] <= 16'h0000;
      coeffs_in_data_log_force[6426] <= 16'h0000;
      coeffs_in_data_log_force[6427] <= 16'h0000;
      coeffs_in_data_log_force[6428] <= 16'h0000;
      coeffs_in_data_log_force[6429] <= 16'h0000;
      coeffs_in_data_log_force[6430] <= 16'h0000;
      coeffs_in_data_log_force[6431] <= 16'h0000;
      coeffs_in_data_log_force[6432] <= 16'h0000;
      coeffs_in_data_log_force[6433] <= 16'h0000;
      coeffs_in_data_log_force[6434] <= 16'h0000;
      coeffs_in_data_log_force[6435] <= 16'h0000;
      coeffs_in_data_log_force[6436] <= 16'h0000;
      coeffs_in_data_log_force[6437] <= 16'h0000;
      coeffs_in_data_log_force[6438] <= 16'h0000;
      coeffs_in_data_log_force[6439] <= 16'h0000;
      coeffs_in_data_log_force[6440] <= 16'h0000;
      coeffs_in_data_log_force[6441] <= 16'h0000;
      coeffs_in_data_log_force[6442] <= 16'h0000;
      coeffs_in_data_log_force[6443] <= 16'h0000;
      coeffs_in_data_log_force[6444] <= 16'h0000;
      coeffs_in_data_log_force[6445] <= 16'h0000;
      coeffs_in_data_log_force[6446] <= 16'h0000;
      coeffs_in_data_log_force[6447] <= 16'h0000;
      coeffs_in_data_log_force[6448] <= 16'h0000;
      coeffs_in_data_log_force[6449] <= 16'h0000;
      coeffs_in_data_log_force[6450] <= 16'h0000;
      coeffs_in_data_log_force[6451] <= 16'h0000;
      coeffs_in_data_log_force[6452] <= 16'h0000;
      coeffs_in_data_log_force[6453] <= 16'h0000;
      coeffs_in_data_log_force[6454] <= 16'h0000;
      coeffs_in_data_log_force[6455] <= 16'h0000;
      coeffs_in_data_log_force[6456] <= 16'h0000;
      coeffs_in_data_log_force[6457] <= 16'h0000;
      coeffs_in_data_log_force[6458] <= 16'h0000;
      coeffs_in_data_log_force[6459] <= 16'h0000;
      coeffs_in_data_log_force[6460] <= 16'h0000;
      coeffs_in_data_log_force[6461] <= 16'h0000;
      coeffs_in_data_log_force[6462] <= 16'h0000;
      coeffs_in_data_log_force[6463] <= 16'h0000;
      coeffs_in_data_log_force[6464] <= 16'h0000;
      coeffs_in_data_log_force[6465] <= 16'h0000;
      coeffs_in_data_log_force[6466] <= 16'h0000;
      coeffs_in_data_log_force[6467] <= 16'h0000;
      coeffs_in_data_log_force[6468] <= 16'h0000;
      coeffs_in_data_log_force[6469] <= 16'h0000;
      coeffs_in_data_log_force[6470] <= 16'h0000;
      coeffs_in_data_log_force[6471] <= 16'h0000;
      coeffs_in_data_log_force[6472] <= 16'h0000;
      coeffs_in_data_log_force[6473] <= 16'h0000;
      coeffs_in_data_log_force[6474] <= 16'h0000;
      coeffs_in_data_log_force[6475] <= 16'h0000;
      coeffs_in_data_log_force[6476] <= 16'h0000;
      coeffs_in_data_log_force[6477] <= 16'h0000;
      coeffs_in_data_log_force[6478] <= 16'h0000;
      coeffs_in_data_log_force[6479] <= 16'h0000;
      coeffs_in_data_log_force[6480] <= 16'h0000;
      coeffs_in_data_log_force[6481] <= 16'h0000;
      coeffs_in_data_log_force[6482] <= 16'h0000;
      coeffs_in_data_log_force[6483] <= 16'h0000;
      coeffs_in_data_log_force[6484] <= 16'h0000;
      coeffs_in_data_log_force[6485] <= 16'h0000;
      coeffs_in_data_log_force[6486] <= 16'h0000;
      coeffs_in_data_log_force[6487] <= 16'h0000;
      coeffs_in_data_log_force[6488] <= 16'h0000;
      coeffs_in_data_log_force[6489] <= 16'h0000;
      coeffs_in_data_log_force[6490] <= 16'h0000;
      coeffs_in_data_log_force[6491] <= 16'h0000;
      coeffs_in_data_log_force[6492] <= 16'h0000;
      coeffs_in_data_log_force[6493] <= 16'h0000;
      coeffs_in_data_log_force[6494] <= 16'h0000;
      coeffs_in_data_log_force[6495] <= 16'h0000;
      coeffs_in_data_log_force[6496] <= 16'h0000;
      coeffs_in_data_log_force[6497] <= 16'h0000;
      coeffs_in_data_log_force[6498] <= 16'h0000;
      coeffs_in_data_log_force[6499] <= 16'h0000;
      coeffs_in_data_log_force[6500] <= 16'h0000;
      coeffs_in_data_log_force[6501] <= 16'h0000;
      coeffs_in_data_log_force[6502] <= 16'h0000;
      coeffs_in_data_log_force[6503] <= 16'h0000;
      coeffs_in_data_log_force[6504] <= 16'h0000;
      coeffs_in_data_log_force[6505] <= 16'h0000;
      coeffs_in_data_log_force[6506] <= 16'h0000;
      coeffs_in_data_log_force[6507] <= 16'h0000;
      coeffs_in_data_log_force[6508] <= 16'h0000;
      coeffs_in_data_log_force[6509] <= 16'h0000;
      coeffs_in_data_log_force[6510] <= 16'h0000;
      coeffs_in_data_log_force[6511] <= 16'h0000;
      coeffs_in_data_log_force[6512] <= 16'h0000;
      coeffs_in_data_log_force[6513] <= 16'h0000;
      coeffs_in_data_log_force[6514] <= 16'h0000;
      coeffs_in_data_log_force[6515] <= 16'h0000;
      coeffs_in_data_log_force[6516] <= 16'h0000;
      coeffs_in_data_log_force[6517] <= 16'h0000;
      coeffs_in_data_log_force[6518] <= 16'h0000;
      coeffs_in_data_log_force[6519] <= 16'h0000;
      coeffs_in_data_log_force[6520] <= 16'h0000;
      coeffs_in_data_log_force[6521] <= 16'h0000;
      coeffs_in_data_log_force[6522] <= 16'h0000;
      coeffs_in_data_log_force[6523] <= 16'h0000;
      coeffs_in_data_log_force[6524] <= 16'h0000;
      coeffs_in_data_log_force[6525] <= 16'h0000;
      coeffs_in_data_log_force[6526] <= 16'h0000;
      coeffs_in_data_log_force[6527] <= 16'h0000;
      coeffs_in_data_log_force[6528] <= 16'h0000;
      coeffs_in_data_log_force[6529] <= 16'h0000;
      coeffs_in_data_log_force[6530] <= 16'h0000;
      coeffs_in_data_log_force[6531] <= 16'h0000;
      coeffs_in_data_log_force[6532] <= 16'h0000;
      coeffs_in_data_log_force[6533] <= 16'h0000;
      coeffs_in_data_log_force[6534] <= 16'h0000;
      coeffs_in_data_log_force[6535] <= 16'h0000;
      coeffs_in_data_log_force[6536] <= 16'h0000;
      coeffs_in_data_log_force[6537] <= 16'h0000;
      coeffs_in_data_log_force[6538] <= 16'h0000;
      coeffs_in_data_log_force[6539] <= 16'h0000;
      coeffs_in_data_log_force[6540] <= 16'h0000;
      coeffs_in_data_log_force[6541] <= 16'h0000;
      coeffs_in_data_log_force[6542] <= 16'h0000;
      coeffs_in_data_log_force[6543] <= 16'h0000;
      coeffs_in_data_log_force[6544] <= 16'h0000;
      coeffs_in_data_log_force[6545] <= 16'h0000;
      coeffs_in_data_log_force[6546] <= 16'h0000;
      coeffs_in_data_log_force[6547] <= 16'h0000;
      coeffs_in_data_log_force[6548] <= 16'h0000;
      coeffs_in_data_log_force[6549] <= 16'h0000;
      coeffs_in_data_log_force[6550] <= 16'h0000;
      coeffs_in_data_log_force[6551] <= 16'h0000;
      coeffs_in_data_log_force[6552] <= 16'h0000;
      coeffs_in_data_log_force[6553] <= 16'h0000;
      coeffs_in_data_log_force[6554] <= 16'h0000;
      coeffs_in_data_log_force[6555] <= 16'h0000;
      coeffs_in_data_log_force[6556] <= 16'h0000;
      coeffs_in_data_log_force[6557] <= 16'h0000;
      coeffs_in_data_log_force[6558] <= 16'h0000;
      coeffs_in_data_log_force[6559] <= 16'h0000;
      coeffs_in_data_log_force[6560] <= 16'h0000;
      coeffs_in_data_log_force[6561] <= 16'h0000;
      coeffs_in_data_log_force[6562] <= 16'h0000;
      coeffs_in_data_log_force[6563] <= 16'h0000;
      coeffs_in_data_log_force[6564] <= 16'h0000;
      coeffs_in_data_log_force[6565] <= 16'h0000;
      coeffs_in_data_log_force[6566] <= 16'h0000;
      coeffs_in_data_log_force[6567] <= 16'h0000;
      coeffs_in_data_log_force[6568] <= 16'h0000;
      coeffs_in_data_log_force[6569] <= 16'h0000;
      coeffs_in_data_log_force[6570] <= 16'h0000;
      coeffs_in_data_log_force[6571] <= 16'h0000;
      coeffs_in_data_log_force[6572] <= 16'h0000;
      coeffs_in_data_log_force[6573] <= 16'h0000;
      coeffs_in_data_log_force[6574] <= 16'h0000;
      coeffs_in_data_log_force[6575] <= 16'h0000;
      coeffs_in_data_log_force[6576] <= 16'h0000;
      coeffs_in_data_log_force[6577] <= 16'h0000;
      coeffs_in_data_log_force[6578] <= 16'h0000;
      coeffs_in_data_log_force[6579] <= 16'h0000;
      coeffs_in_data_log_force[6580] <= 16'h0000;
      coeffs_in_data_log_force[6581] <= 16'h0000;
      coeffs_in_data_log_force[6582] <= 16'h0000;
      coeffs_in_data_log_force[6583] <= 16'h0000;
      coeffs_in_data_log_force[6584] <= 16'h0000;
      coeffs_in_data_log_force[6585] <= 16'h0000;
      coeffs_in_data_log_force[6586] <= 16'h0000;
      coeffs_in_data_log_force[6587] <= 16'h0000;
      coeffs_in_data_log_force[6588] <= 16'h0000;
      coeffs_in_data_log_force[6589] <= 16'h0000;
      coeffs_in_data_log_force[6590] <= 16'h0000;
      coeffs_in_data_log_force[6591] <= 16'h0000;
      coeffs_in_data_log_force[6592] <= 16'h0000;
      coeffs_in_data_log_force[6593] <= 16'h0000;
      coeffs_in_data_log_force[6594] <= 16'h0000;
      coeffs_in_data_log_force[6595] <= 16'h0000;
      coeffs_in_data_log_force[6596] <= 16'h0000;
      coeffs_in_data_log_force[6597] <= 16'h0000;
      coeffs_in_data_log_force[6598] <= 16'h0000;
      coeffs_in_data_log_force[6599] <= 16'h0000;
      coeffs_in_data_log_force[6600] <= 16'h0000;
      coeffs_in_data_log_force[6601] <= 16'h0000;
      coeffs_in_data_log_force[6602] <= 16'h0000;
      coeffs_in_data_log_force[6603] <= 16'h0000;
      coeffs_in_data_log_force[6604] <= 16'h0000;
      coeffs_in_data_log_force[6605] <= 16'h0000;
      coeffs_in_data_log_force[6606] <= 16'h0000;
      coeffs_in_data_log_force[6607] <= 16'h0000;
      coeffs_in_data_log_force[6608] <= 16'h0000;
      coeffs_in_data_log_force[6609] <= 16'h0000;
      coeffs_in_data_log_force[6610] <= 16'h0000;
      coeffs_in_data_log_force[6611] <= 16'h0000;
      coeffs_in_data_log_force[6612] <= 16'h0000;
      coeffs_in_data_log_force[6613] <= 16'h0000;
      coeffs_in_data_log_force[6614] <= 16'h0000;
      coeffs_in_data_log_force[6615] <= 16'h0000;
      coeffs_in_data_log_force[6616] <= 16'h0000;
      coeffs_in_data_log_force[6617] <= 16'h0000;
      coeffs_in_data_log_force[6618] <= 16'h0000;
      coeffs_in_data_log_force[6619] <= 16'h0000;
      coeffs_in_data_log_force[6620] <= 16'h0000;
      coeffs_in_data_log_force[6621] <= 16'h0000;
      coeffs_in_data_log_force[6622] <= 16'h0000;
      coeffs_in_data_log_force[6623] <= 16'h0000;
      coeffs_in_data_log_force[6624] <= 16'h0000;
      coeffs_in_data_log_force[6625] <= 16'h0000;
      coeffs_in_data_log_force[6626] <= 16'h0000;
      coeffs_in_data_log_force[6627] <= 16'h0000;
      coeffs_in_data_log_force[6628] <= 16'h0000;
      coeffs_in_data_log_force[6629] <= 16'h0000;
      coeffs_in_data_log_force[6630] <= 16'h0000;
      coeffs_in_data_log_force[6631] <= 16'h0000;
      coeffs_in_data_log_force[6632] <= 16'h0000;
      coeffs_in_data_log_force[6633] <= 16'h0000;
      coeffs_in_data_log_force[6634] <= 16'h0000;
      coeffs_in_data_log_force[6635] <= 16'h0000;
      coeffs_in_data_log_force[6636] <= 16'h0000;
      coeffs_in_data_log_force[6637] <= 16'h0000;
      coeffs_in_data_log_force[6638] <= 16'h0000;
      coeffs_in_data_log_force[6639] <= 16'h0000;
      coeffs_in_data_log_force[6640] <= 16'h0000;
      coeffs_in_data_log_force[6641] <= 16'h0000;
      coeffs_in_data_log_force[6642] <= 16'h0000;
      coeffs_in_data_log_force[6643] <= 16'h0000;
      coeffs_in_data_log_force[6644] <= 16'h0000;
      coeffs_in_data_log_force[6645] <= 16'h0000;
      coeffs_in_data_log_force[6646] <= 16'h0000;
      coeffs_in_data_log_force[6647] <= 16'h0000;
      coeffs_in_data_log_force[6648] <= 16'h0000;
      coeffs_in_data_log_force[6649] <= 16'h0000;
      coeffs_in_data_log_force[6650] <= 16'h0000;
      coeffs_in_data_log_force[6651] <= 16'h0000;
      coeffs_in_data_log_force[6652] <= 16'h0000;
      coeffs_in_data_log_force[6653] <= 16'h0000;
      coeffs_in_data_log_force[6654] <= 16'h0000;
      coeffs_in_data_log_force[6655] <= 16'h0000;
      coeffs_in_data_log_force[6656] <= 16'h0000;
      coeffs_in_data_log_force[6657] <= 16'h0000;
      coeffs_in_data_log_force[6658] <= 16'h0000;
      coeffs_in_data_log_force[6659] <= 16'h0000;
      coeffs_in_data_log_force[6660] <= 16'h0000;
      coeffs_in_data_log_force[6661] <= 16'h0000;
      coeffs_in_data_log_force[6662] <= 16'h0000;
      coeffs_in_data_log_force[6663] <= 16'h0000;
      coeffs_in_data_log_force[6664] <= 16'h0000;
      coeffs_in_data_log_force[6665] <= 16'h0000;
      coeffs_in_data_log_force[6666] <= 16'h0000;
      coeffs_in_data_log_force[6667] <= 16'h0000;
      coeffs_in_data_log_force[6668] <= 16'h0000;
      coeffs_in_data_log_force[6669] <= 16'h0000;
      coeffs_in_data_log_force[6670] <= 16'h0000;
      coeffs_in_data_log_force[6671] <= 16'h0000;
      coeffs_in_data_log_force[6672] <= 16'h0000;
      coeffs_in_data_log_force[6673] <= 16'h0000;
      coeffs_in_data_log_force[6674] <= 16'h0000;
      coeffs_in_data_log_force[6675] <= 16'h0000;
      coeffs_in_data_log_force[6676] <= 16'h0000;
      coeffs_in_data_log_force[6677] <= 16'h0000;
      coeffs_in_data_log_force[6678] <= 16'h0000;
      coeffs_in_data_log_force[6679] <= 16'h0000;
      coeffs_in_data_log_force[6680] <= 16'h0000;
      coeffs_in_data_log_force[6681] <= 16'h0000;
      coeffs_in_data_log_force[6682] <= 16'h0000;
      coeffs_in_data_log_force[6683] <= 16'h0000;
      coeffs_in_data_log_force[6684] <= 16'h0000;
      coeffs_in_data_log_force[6685] <= 16'h0000;
      coeffs_in_data_log_force[6686] <= 16'h0000;
      coeffs_in_data_log_force[6687] <= 16'h0000;
      coeffs_in_data_log_force[6688] <= 16'h0000;
      coeffs_in_data_log_force[6689] <= 16'h0000;
      coeffs_in_data_log_force[6690] <= 16'h0000;
      coeffs_in_data_log_force[6691] <= 16'h0000;
      coeffs_in_data_log_force[6692] <= 16'h0000;
      coeffs_in_data_log_force[6693] <= 16'h0000;
      coeffs_in_data_log_force[6694] <= 16'h0000;
      coeffs_in_data_log_force[6695] <= 16'h0000;
      coeffs_in_data_log_force[6696] <= 16'h0000;
      coeffs_in_data_log_force[6697] <= 16'h0000;
      coeffs_in_data_log_force[6698] <= 16'h0000;
      coeffs_in_data_log_force[6699] <= 16'h0000;
      coeffs_in_data_log_force[6700] <= 16'h0000;
      coeffs_in_data_log_force[6701] <= 16'h0000;
      coeffs_in_data_log_force[6702] <= 16'h0000;
      coeffs_in_data_log_force[6703] <= 16'h0000;
      coeffs_in_data_log_force[6704] <= 16'h0000;
      coeffs_in_data_log_force[6705] <= 16'h0000;
      coeffs_in_data_log_force[6706] <= 16'h0000;
      coeffs_in_data_log_force[6707] <= 16'h0000;
      coeffs_in_data_log_force[6708] <= 16'h0000;
      coeffs_in_data_log_force[6709] <= 16'h0000;
      coeffs_in_data_log_force[6710] <= 16'h0000;
      coeffs_in_data_log_force[6711] <= 16'h0000;
      coeffs_in_data_log_force[6712] <= 16'h0000;
      coeffs_in_data_log_force[6713] <= 16'h0000;
      coeffs_in_data_log_force[6714] <= 16'h0000;
      coeffs_in_data_log_force[6715] <= 16'h0000;
      coeffs_in_data_log_force[6716] <= 16'h0000;
      coeffs_in_data_log_force[6717] <= 16'h0000;
      coeffs_in_data_log_force[6718] <= 16'h0000;
      coeffs_in_data_log_force[6719] <= 16'h0000;
      coeffs_in_data_log_force[6720] <= 16'h0000;
      coeffs_in_data_log_force[6721] <= 16'h0000;
      coeffs_in_data_log_force[6722] <= 16'h0000;
      coeffs_in_data_log_force[6723] <= 16'h0000;
      coeffs_in_data_log_force[6724] <= 16'h0000;
      coeffs_in_data_log_force[6725] <= 16'h0000;
      coeffs_in_data_log_force[6726] <= 16'h0000;
      coeffs_in_data_log_force[6727] <= 16'h0000;
      coeffs_in_data_log_force[6728] <= 16'h0000;
      coeffs_in_data_log_force[6729] <= 16'h0000;
      coeffs_in_data_log_force[6730] <= 16'h0000;
      coeffs_in_data_log_force[6731] <= 16'h0000;
      coeffs_in_data_log_force[6732] <= 16'h0000;
      coeffs_in_data_log_force[6733] <= 16'h0000;
      coeffs_in_data_log_force[6734] <= 16'h0000;
      coeffs_in_data_log_force[6735] <= 16'h0000;
      coeffs_in_data_log_force[6736] <= 16'h0000;
      coeffs_in_data_log_force[6737] <= 16'h0000;
      coeffs_in_data_log_force[6738] <= 16'h0000;
      coeffs_in_data_log_force[6739] <= 16'h0000;
      coeffs_in_data_log_force[6740] <= 16'h0000;
      coeffs_in_data_log_force[6741] <= 16'h0000;
      coeffs_in_data_log_force[6742] <= 16'h0000;
      coeffs_in_data_log_force[6743] <= 16'h0000;
      coeffs_in_data_log_force[6744] <= 16'h0000;
      coeffs_in_data_log_force[6745] <= 16'h0000;
      coeffs_in_data_log_force[6746] <= 16'h0000;
      coeffs_in_data_log_force[6747] <= 16'h0000;
      coeffs_in_data_log_force[6748] <= 16'h0000;
      coeffs_in_data_log_force[6749] <= 16'h0000;
      coeffs_in_data_log_force[6750] <= 16'h0000;
      coeffs_in_data_log_force[6751] <= 16'h0000;
      coeffs_in_data_log_force[6752] <= 16'h0000;
      coeffs_in_data_log_force[6753] <= 16'h0000;
      coeffs_in_data_log_force[6754] <= 16'h0000;
      coeffs_in_data_log_force[6755] <= 16'h0000;
      coeffs_in_data_log_force[6756] <= 16'h0000;
      coeffs_in_data_log_force[6757] <= 16'h0000;
      coeffs_in_data_log_force[6758] <= 16'h0000;
      coeffs_in_data_log_force[6759] <= 16'h0000;
      coeffs_in_data_log_force[6760] <= 16'h0000;
      coeffs_in_data_log_force[6761] <= 16'h0000;
      coeffs_in_data_log_force[6762] <= 16'h0000;
      coeffs_in_data_log_force[6763] <= 16'h0000;
      coeffs_in_data_log_force[6764] <= 16'h0000;
      coeffs_in_data_log_force[6765] <= 16'h0000;
      coeffs_in_data_log_force[6766] <= 16'h0000;
      coeffs_in_data_log_force[6767] <= 16'h0000;
      coeffs_in_data_log_force[6768] <= 16'h0000;
      coeffs_in_data_log_force[6769] <= 16'h0000;
      coeffs_in_data_log_force[6770] <= 16'h0000;
      coeffs_in_data_log_force[6771] <= 16'h0000;
      coeffs_in_data_log_force[6772] <= 16'h0000;
      coeffs_in_data_log_force[6773] <= 16'h0000;
      coeffs_in_data_log_force[6774] <= 16'h0000;
      coeffs_in_data_log_force[6775] <= 16'h0000;
      coeffs_in_data_log_force[6776] <= 16'h0000;
      coeffs_in_data_log_force[6777] <= 16'h0000;
      coeffs_in_data_log_force[6778] <= 16'h0000;
      coeffs_in_data_log_force[6779] <= 16'h0000;
      coeffs_in_data_log_force[6780] <= 16'h0000;
      coeffs_in_data_log_force[6781] <= 16'h0000;
      coeffs_in_data_log_force[6782] <= 16'h0000;
      coeffs_in_data_log_force[6783] <= 16'h0000;
      coeffs_in_data_log_force[6784] <= 16'h0000;
      coeffs_in_data_log_force[6785] <= 16'h0000;
      coeffs_in_data_log_force[6786] <= 16'h0000;
      coeffs_in_data_log_force[6787] <= 16'h0000;
      coeffs_in_data_log_force[6788] <= 16'h0000;
      coeffs_in_data_log_force[6789] <= 16'h0000;
      coeffs_in_data_log_force[6790] <= 16'h0000;
      coeffs_in_data_log_force[6791] <= 16'h0000;
      coeffs_in_data_log_force[6792] <= 16'h0000;
      coeffs_in_data_log_force[6793] <= 16'h0000;
      coeffs_in_data_log_force[6794] <= 16'h0000;
      coeffs_in_data_log_force[6795] <= 16'h0000;
      coeffs_in_data_log_force[6796] <= 16'h0000;
      coeffs_in_data_log_force[6797] <= 16'h0000;
      coeffs_in_data_log_force[6798] <= 16'h0000;
      coeffs_in_data_log_force[6799] <= 16'h0000;
      coeffs_in_data_log_force[6800] <= 16'h0000;
      coeffs_in_data_log_force[6801] <= 16'h0000;
      coeffs_in_data_log_force[6802] <= 16'h0000;
      coeffs_in_data_log_force[6803] <= 16'h0000;
      coeffs_in_data_log_force[6804] <= 16'h0000;
      coeffs_in_data_log_force[6805] <= 16'h0000;
      coeffs_in_data_log_force[6806] <= 16'h0000;
      coeffs_in_data_log_force[6807] <= 16'h0000;
      coeffs_in_data_log_force[6808] <= 16'h0000;
      coeffs_in_data_log_force[6809] <= 16'h0000;
      coeffs_in_data_log_force[6810] <= 16'h0000;
      coeffs_in_data_log_force[6811] <= 16'h0000;
      coeffs_in_data_log_force[6812] <= 16'h0000;
      coeffs_in_data_log_force[6813] <= 16'h0000;
      coeffs_in_data_log_force[6814] <= 16'h0000;
      coeffs_in_data_log_force[6815] <= 16'h0000;
      coeffs_in_data_log_force[6816] <= 16'h0000;
      coeffs_in_data_log_force[6817] <= 16'h0000;
      coeffs_in_data_log_force[6818] <= 16'h0000;
      coeffs_in_data_log_force[6819] <= 16'h0000;
      coeffs_in_data_log_force[6820] <= 16'h0000;
      coeffs_in_data_log_force[6821] <= 16'h0000;
      coeffs_in_data_log_force[6822] <= 16'h0000;
      coeffs_in_data_log_force[6823] <= 16'h0000;
      coeffs_in_data_log_force[6824] <= 16'h0000;
      coeffs_in_data_log_force[6825] <= 16'h0000;
      coeffs_in_data_log_force[6826] <= 16'h0000;
      coeffs_in_data_log_force[6827] <= 16'h0000;
      coeffs_in_data_log_force[6828] <= 16'h0000;
      coeffs_in_data_log_force[6829] <= 16'h0000;
      coeffs_in_data_log_force[6830] <= 16'h0000;
      coeffs_in_data_log_force[6831] <= 16'h0000;
      coeffs_in_data_log_force[6832] <= 16'h0000;
      coeffs_in_data_log_force[6833] <= 16'h0000;
      coeffs_in_data_log_force[6834] <= 16'h0000;
      coeffs_in_data_log_force[6835] <= 16'h0000;
      coeffs_in_data_log_force[6836] <= 16'h0000;
      coeffs_in_data_log_force[6837] <= 16'h0000;
      coeffs_in_data_log_force[6838] <= 16'h0000;
      coeffs_in_data_log_force[6839] <= 16'h0000;
      coeffs_in_data_log_force[6840] <= 16'h0000;
      coeffs_in_data_log_force[6841] <= 16'h0000;
      coeffs_in_data_log_force[6842] <= 16'h0000;
      coeffs_in_data_log_force[6843] <= 16'h0000;
      coeffs_in_data_log_force[6844] <= 16'h0000;
      coeffs_in_data_log_force[6845] <= 16'h0000;
      coeffs_in_data_log_force[6846] <= 16'h0000;
      coeffs_in_data_log_force[6847] <= 16'h0000;
      coeffs_in_data_log_force[6848] <= 16'h0000;
      coeffs_in_data_log_force[6849] <= 16'h0000;
      coeffs_in_data_log_force[6850] <= 16'h0000;
      coeffs_in_data_log_force[6851] <= 16'h0000;
      coeffs_in_data_log_force[6852] <= 16'h0000;
      coeffs_in_data_log_force[6853] <= 16'h0000;
      coeffs_in_data_log_force[6854] <= 16'h0000;
      coeffs_in_data_log_force[6855] <= 16'h0000;
      coeffs_in_data_log_force[6856] <= 16'h0000;
      coeffs_in_data_log_force[6857] <= 16'h0000;
      coeffs_in_data_log_force[6858] <= 16'h0000;
      coeffs_in_data_log_force[6859] <= 16'h0000;
      coeffs_in_data_log_force[6860] <= 16'h0000;
      coeffs_in_data_log_force[6861] <= 16'h0000;
      coeffs_in_data_log_force[6862] <= 16'h0000;
      coeffs_in_data_log_force[6863] <= 16'h0000;
      coeffs_in_data_log_force[6864] <= 16'h0000;
      coeffs_in_data_log_force[6865] <= 16'h0000;
      coeffs_in_data_log_force[6866] <= 16'h0000;
      coeffs_in_data_log_force[6867] <= 16'h0000;
      coeffs_in_data_log_force[6868] <= 16'h0000;
      coeffs_in_data_log_force[6869] <= 16'h0000;
      coeffs_in_data_log_force[6870] <= 16'h0000;
      coeffs_in_data_log_force[6871] <= 16'h0000;
      coeffs_in_data_log_force[6872] <= 16'h0000;
      coeffs_in_data_log_force[6873] <= 16'h0000;
      coeffs_in_data_log_force[6874] <= 16'h0000;
      coeffs_in_data_log_force[6875] <= 16'h0000;
      coeffs_in_data_log_force[6876] <= 16'h0000;
      coeffs_in_data_log_force[6877] <= 16'h0000;
      coeffs_in_data_log_force[6878] <= 16'h0000;
      coeffs_in_data_log_force[6879] <= 16'h0000;
      coeffs_in_data_log_force[6880] <= 16'h0000;
      coeffs_in_data_log_force[6881] <= 16'h0000;
      coeffs_in_data_log_force[6882] <= 16'h0000;
      coeffs_in_data_log_force[6883] <= 16'h0000;
      coeffs_in_data_log_force[6884] <= 16'h0000;
      coeffs_in_data_log_force[6885] <= 16'h0000;
      coeffs_in_data_log_force[6886] <= 16'h0000;
      coeffs_in_data_log_force[6887] <= 16'h0000;
      coeffs_in_data_log_force[6888] <= 16'h0000;
      coeffs_in_data_log_force[6889] <= 16'h0000;
      coeffs_in_data_log_force[6890] <= 16'h0000;
      coeffs_in_data_log_force[6891] <= 16'h0000;
      coeffs_in_data_log_force[6892] <= 16'h0000;
      coeffs_in_data_log_force[6893] <= 16'h0000;
      coeffs_in_data_log_force[6894] <= 16'h0000;
      coeffs_in_data_log_force[6895] <= 16'h0000;
      coeffs_in_data_log_force[6896] <= 16'h0000;
      coeffs_in_data_log_force[6897] <= 16'h0000;
      coeffs_in_data_log_force[6898] <= 16'h0000;
      coeffs_in_data_log_force[6899] <= 16'h0000;
      coeffs_in_data_log_force[6900] <= 16'h0000;
      coeffs_in_data_log_force[6901] <= 16'h0000;
      coeffs_in_data_log_force[6902] <= 16'h0000;
      coeffs_in_data_log_force[6903] <= 16'h0000;
      coeffs_in_data_log_force[6904] <= 16'h0000;
      coeffs_in_data_log_force[6905] <= 16'h0000;
      coeffs_in_data_log_force[6906] <= 16'h0000;
      coeffs_in_data_log_force[6907] <= 16'h0000;
      coeffs_in_data_log_force[6908] <= 16'h0000;
      coeffs_in_data_log_force[6909] <= 16'h0000;
      coeffs_in_data_log_force[6910] <= 16'h0000;
      coeffs_in_data_log_force[6911] <= 16'h0000;
      coeffs_in_data_log_force[6912] <= 16'h0000;
      coeffs_in_data_log_force[6913] <= 16'h0000;
      coeffs_in_data_log_force[6914] <= 16'h0000;
      coeffs_in_data_log_force[6915] <= 16'h0000;
      coeffs_in_data_log_force[6916] <= 16'h0000;
      coeffs_in_data_log_force[6917] <= 16'h0000;
      coeffs_in_data_log_force[6918] <= 16'h0000;
      coeffs_in_data_log_force[6919] <= 16'h0000;
      coeffs_in_data_log_force[6920] <= 16'h0000;
      coeffs_in_data_log_force[6921] <= 16'h0000;
      coeffs_in_data_log_force[6922] <= 16'h0000;
      coeffs_in_data_log_force[6923] <= 16'h0000;
      coeffs_in_data_log_force[6924] <= 16'h0000;
      coeffs_in_data_log_force[6925] <= 16'h0000;
      coeffs_in_data_log_force[6926] <= 16'h0000;
      coeffs_in_data_log_force[6927] <= 16'h0000;
      coeffs_in_data_log_force[6928] <= 16'h0000;
      coeffs_in_data_log_force[6929] <= 16'h0000;
      coeffs_in_data_log_force[6930] <= 16'h0000;
      coeffs_in_data_log_force[6931] <= 16'h0000;
      coeffs_in_data_log_force[6932] <= 16'h0000;
      coeffs_in_data_log_force[6933] <= 16'h0000;
      coeffs_in_data_log_force[6934] <= 16'h0000;
      coeffs_in_data_log_force[6935] <= 16'h0000;
      coeffs_in_data_log_force[6936] <= 16'h0000;
      coeffs_in_data_log_force[6937] <= 16'h0000;
      coeffs_in_data_log_force[6938] <= 16'h0000;
      coeffs_in_data_log_force[6939] <= 16'h0000;
      coeffs_in_data_log_force[6940] <= 16'h0000;
      coeffs_in_data_log_force[6941] <= 16'h0000;
      coeffs_in_data_log_force[6942] <= 16'h0000;
      coeffs_in_data_log_force[6943] <= 16'h0000;
      coeffs_in_data_log_force[6944] <= 16'h0000;
      coeffs_in_data_log_force[6945] <= 16'h0000;
      coeffs_in_data_log_force[6946] <= 16'h0000;
      coeffs_in_data_log_force[6947] <= 16'h0000;
      coeffs_in_data_log_force[6948] <= 16'h0000;
      coeffs_in_data_log_force[6949] <= 16'h0000;
      coeffs_in_data_log_force[6950] <= 16'h0000;
      coeffs_in_data_log_force[6951] <= 16'h0000;
      coeffs_in_data_log_force[6952] <= 16'h0000;
      coeffs_in_data_log_force[6953] <= 16'h0000;
      coeffs_in_data_log_force[6954] <= 16'h0000;
      coeffs_in_data_log_force[6955] <= 16'h0000;
      coeffs_in_data_log_force[6956] <= 16'h0000;
      coeffs_in_data_log_force[6957] <= 16'h0000;
      coeffs_in_data_log_force[6958] <= 16'h0000;
      coeffs_in_data_log_force[6959] <= 16'h0000;
      coeffs_in_data_log_force[6960] <= 16'h0000;
      coeffs_in_data_log_force[6961] <= 16'h0000;
      coeffs_in_data_log_force[6962] <= 16'h0000;
      coeffs_in_data_log_force[6963] <= 16'h0000;
      coeffs_in_data_log_force[6964] <= 16'h0000;
      coeffs_in_data_log_force[6965] <= 16'h0000;
      coeffs_in_data_log_force[6966] <= 16'h0000;
      coeffs_in_data_log_force[6967] <= 16'h0000;
      coeffs_in_data_log_force[6968] <= 16'h0000;
      coeffs_in_data_log_force[6969] <= 16'h0000;
      coeffs_in_data_log_force[6970] <= 16'h0000;
      coeffs_in_data_log_force[6971] <= 16'h0000;
      coeffs_in_data_log_force[6972] <= 16'h0000;
      coeffs_in_data_log_force[6973] <= 16'h0000;
      coeffs_in_data_log_force[6974] <= 16'h0000;
      coeffs_in_data_log_force[6975] <= 16'h0000;
      coeffs_in_data_log_force[6976] <= 16'h0000;
      coeffs_in_data_log_force[6977] <= 16'h0000;
      coeffs_in_data_log_force[6978] <= 16'h0000;
      coeffs_in_data_log_force[6979] <= 16'h0000;
      coeffs_in_data_log_force[6980] <= 16'h0000;
      coeffs_in_data_log_force[6981] <= 16'h0000;
      coeffs_in_data_log_force[6982] <= 16'h0000;
      coeffs_in_data_log_force[6983] <= 16'h0000;
      coeffs_in_data_log_force[6984] <= 16'h0000;
      coeffs_in_data_log_force[6985] <= 16'h0000;
      coeffs_in_data_log_force[6986] <= 16'h0000;
      coeffs_in_data_log_force[6987] <= 16'h0000;
      coeffs_in_data_log_force[6988] <= 16'h0000;
      coeffs_in_data_log_force[6989] <= 16'h0000;
      coeffs_in_data_log_force[6990] <= 16'h0000;
      coeffs_in_data_log_force[6991] <= 16'h0000;
      coeffs_in_data_log_force[6992] <= 16'h0000;
      coeffs_in_data_log_force[6993] <= 16'h0000;
      coeffs_in_data_log_force[6994] <= 16'h0000;
      coeffs_in_data_log_force[6995] <= 16'h0000;
      coeffs_in_data_log_force[6996] <= 16'h0000;
      coeffs_in_data_log_force[6997] <= 16'h0000;
      coeffs_in_data_log_force[6998] <= 16'h0000;
      coeffs_in_data_log_force[6999] <= 16'h0000;
      coeffs_in_data_log_force[7000] <= 16'h0000;
      coeffs_in_data_log_force[7001] <= 16'h0000;
      coeffs_in_data_log_force[7002] <= 16'h0000;
      coeffs_in_data_log_force[7003] <= 16'h0000;
      coeffs_in_data_log_force[7004] <= 16'h0000;
      coeffs_in_data_log_force[7005] <= 16'h0000;
      coeffs_in_data_log_force[7006] <= 16'h0000;
      coeffs_in_data_log_force[7007] <= 16'h0000;
      coeffs_in_data_log_force[7008] <= 16'h0000;
      coeffs_in_data_log_force[7009] <= 16'h0000;
      coeffs_in_data_log_force[7010] <= 16'h0000;
      coeffs_in_data_log_force[7011] <= 16'h0000;
      coeffs_in_data_log_force[7012] <= 16'h0000;
      coeffs_in_data_log_force[7013] <= 16'h0000;
      coeffs_in_data_log_force[7014] <= 16'h0000;
      coeffs_in_data_log_force[7015] <= 16'h0000;
      coeffs_in_data_log_force[7016] <= 16'h0000;
      coeffs_in_data_log_force[7017] <= 16'h0000;
      coeffs_in_data_log_force[7018] <= 16'h0000;
      coeffs_in_data_log_force[7019] <= 16'h0000;
      coeffs_in_data_log_force[7020] <= 16'h0000;
      coeffs_in_data_log_force[7021] <= 16'h0000;
      coeffs_in_data_log_force[7022] <= 16'h0000;
      coeffs_in_data_log_force[7023] <= 16'h0000;
      coeffs_in_data_log_force[7024] <= 16'h0000;
      coeffs_in_data_log_force[7025] <= 16'h0000;
      coeffs_in_data_log_force[7026] <= 16'h0000;
      coeffs_in_data_log_force[7027] <= 16'h0000;
      coeffs_in_data_log_force[7028] <= 16'h0000;
      coeffs_in_data_log_force[7029] <= 16'h0000;
      coeffs_in_data_log_force[7030] <= 16'h0000;
      coeffs_in_data_log_force[7031] <= 16'h0000;
      coeffs_in_data_log_force[7032] <= 16'h0000;
      coeffs_in_data_log_force[7033] <= 16'h0000;
      coeffs_in_data_log_force[7034] <= 16'h0000;
      coeffs_in_data_log_force[7035] <= 16'h0000;
      coeffs_in_data_log_force[7036] <= 16'h0000;
      coeffs_in_data_log_force[7037] <= 16'h0000;
      coeffs_in_data_log_force[7038] <= 16'h0000;
      coeffs_in_data_log_force[7039] <= 16'h0000;
      coeffs_in_data_log_force[7040] <= 16'h0000;
      coeffs_in_data_log_force[7041] <= 16'h0000;
      coeffs_in_data_log_force[7042] <= 16'h0000;
      coeffs_in_data_log_force[7043] <= 16'h0000;
      coeffs_in_data_log_force[7044] <= 16'h0000;
      coeffs_in_data_log_force[7045] <= 16'h0000;
      coeffs_in_data_log_force[7046] <= 16'h0000;
      coeffs_in_data_log_force[7047] <= 16'h0000;
      coeffs_in_data_log_force[7048] <= 16'h0000;
      coeffs_in_data_log_force[7049] <= 16'h0000;
      coeffs_in_data_log_force[7050] <= 16'h0000;
      coeffs_in_data_log_force[7051] <= 16'h0000;
      coeffs_in_data_log_force[7052] <= 16'h0000;
      coeffs_in_data_log_force[7053] <= 16'h0000;
      coeffs_in_data_log_force[7054] <= 16'h0000;
      coeffs_in_data_log_force[7055] <= 16'h0000;
      coeffs_in_data_log_force[7056] <= 16'h0000;
      coeffs_in_data_log_force[7057] <= 16'h0000;
      coeffs_in_data_log_force[7058] <= 16'h0000;
      coeffs_in_data_log_force[7059] <= 16'h0000;
      coeffs_in_data_log_force[7060] <= 16'h0000;
      coeffs_in_data_log_force[7061] <= 16'h0000;
      coeffs_in_data_log_force[7062] <= 16'h0000;
      coeffs_in_data_log_force[7063] <= 16'h0000;
      coeffs_in_data_log_force[7064] <= 16'h0000;
      coeffs_in_data_log_force[7065] <= 16'h0000;
      coeffs_in_data_log_force[7066] <= 16'h0000;
      coeffs_in_data_log_force[7067] <= 16'h0000;
      coeffs_in_data_log_force[7068] <= 16'h0000;
      coeffs_in_data_log_force[7069] <= 16'h0000;
      coeffs_in_data_log_force[7070] <= 16'h0000;
      coeffs_in_data_log_force[7071] <= 16'h0000;
      coeffs_in_data_log_force[7072] <= 16'h0000;
      coeffs_in_data_log_force[7073] <= 16'h0000;
      coeffs_in_data_log_force[7074] <= 16'h0000;
      coeffs_in_data_log_force[7075] <= 16'h0000;
      coeffs_in_data_log_force[7076] <= 16'h0000;
      coeffs_in_data_log_force[7077] <= 16'h0000;
      coeffs_in_data_log_force[7078] <= 16'h0000;
      coeffs_in_data_log_force[7079] <= 16'h0000;
      coeffs_in_data_log_force[7080] <= 16'h0000;
      coeffs_in_data_log_force[7081] <= 16'h0000;
      coeffs_in_data_log_force[7082] <= 16'h0000;
      coeffs_in_data_log_force[7083] <= 16'h0000;
      coeffs_in_data_log_force[7084] <= 16'h0000;
      coeffs_in_data_log_force[7085] <= 16'h0000;
      coeffs_in_data_log_force[7086] <= 16'h0000;
      coeffs_in_data_log_force[7087] <= 16'h0000;
      coeffs_in_data_log_force[7088] <= 16'h0000;
      coeffs_in_data_log_force[7089] <= 16'h0000;
      coeffs_in_data_log_force[7090] <= 16'h0000;
      coeffs_in_data_log_force[7091] <= 16'h0000;
      coeffs_in_data_log_force[7092] <= 16'h0000;
      coeffs_in_data_log_force[7093] <= 16'h0000;
      coeffs_in_data_log_force[7094] <= 16'h0000;
      coeffs_in_data_log_force[7095] <= 16'h0000;
      coeffs_in_data_log_force[7096] <= 16'h0000;
      coeffs_in_data_log_force[7097] <= 16'h0000;
      coeffs_in_data_log_force[7098] <= 16'h0000;
      coeffs_in_data_log_force[7099] <= 16'h0000;
      coeffs_in_data_log_force[7100] <= 16'h0000;
      coeffs_in_data_log_force[7101] <= 16'h0000;
      coeffs_in_data_log_force[7102] <= 16'h0000;
      coeffs_in_data_log_force[7103] <= 16'h0000;
      coeffs_in_data_log_force[7104] <= 16'h0000;
      coeffs_in_data_log_force[7105] <= 16'h0000;
      coeffs_in_data_log_force[7106] <= 16'h0000;
      coeffs_in_data_log_force[7107] <= 16'h0000;
      coeffs_in_data_log_force[7108] <= 16'h0000;
      coeffs_in_data_log_force[7109] <= 16'h0000;
      coeffs_in_data_log_force[7110] <= 16'h0000;
      coeffs_in_data_log_force[7111] <= 16'h0000;
      coeffs_in_data_log_force[7112] <= 16'h0000;
      coeffs_in_data_log_force[7113] <= 16'h0000;
      coeffs_in_data_log_force[7114] <= 16'h0000;
      coeffs_in_data_log_force[7115] <= 16'h0000;
      coeffs_in_data_log_force[7116] <= 16'h0000;
      coeffs_in_data_log_force[7117] <= 16'h0000;
      coeffs_in_data_log_force[7118] <= 16'h0000;
      coeffs_in_data_log_force[7119] <= 16'h0000;
      coeffs_in_data_log_force[7120] <= 16'h0000;
      coeffs_in_data_log_force[7121] <= 16'h0000;
      coeffs_in_data_log_force[7122] <= 16'h0000;
      coeffs_in_data_log_force[7123] <= 16'h0000;
      coeffs_in_data_log_force[7124] <= 16'h0000;
      coeffs_in_data_log_force[7125] <= 16'h0000;
      coeffs_in_data_log_force[7126] <= 16'h0000;
      coeffs_in_data_log_force[7127] <= 16'h0000;
      coeffs_in_data_log_force[7128] <= 16'h0000;
      coeffs_in_data_log_force[7129] <= 16'h0000;
      coeffs_in_data_log_force[7130] <= 16'h0000;
      coeffs_in_data_log_force[7131] <= 16'h0000;
      coeffs_in_data_log_force[7132] <= 16'h0000;
      coeffs_in_data_log_force[7133] <= 16'h0000;
      coeffs_in_data_log_force[7134] <= 16'h0000;
      coeffs_in_data_log_force[7135] <= 16'h0000;
      coeffs_in_data_log_force[7136] <= 16'h0000;
      coeffs_in_data_log_force[7137] <= 16'h0000;
      coeffs_in_data_log_force[7138] <= 16'h0000;
      coeffs_in_data_log_force[7139] <= 16'h0000;
      coeffs_in_data_log_force[7140] <= 16'h0000;
      coeffs_in_data_log_force[7141] <= 16'h0000;
      coeffs_in_data_log_force[7142] <= 16'h0000;
      coeffs_in_data_log_force[7143] <= 16'h0000;
      coeffs_in_data_log_force[7144] <= 16'h0000;
      coeffs_in_data_log_force[7145] <= 16'h0000;
      coeffs_in_data_log_force[7146] <= 16'h0000;
      coeffs_in_data_log_force[7147] <= 16'h0000;
      coeffs_in_data_log_force[7148] <= 16'h0000;
      coeffs_in_data_log_force[7149] <= 16'h0000;
      coeffs_in_data_log_force[7150] <= 16'h0000;
      coeffs_in_data_log_force[7151] <= 16'h0000;
      coeffs_in_data_log_force[7152] <= 16'h0000;
      coeffs_in_data_log_force[7153] <= 16'h0000;
      coeffs_in_data_log_force[7154] <= 16'h0000;
      coeffs_in_data_log_force[7155] <= 16'h0000;
      coeffs_in_data_log_force[7156] <= 16'h0000;
      coeffs_in_data_log_force[7157] <= 16'h0000;
      coeffs_in_data_log_force[7158] <= 16'h0000;
      coeffs_in_data_log_force[7159] <= 16'h0000;
      coeffs_in_data_log_force[7160] <= 16'h0000;
      coeffs_in_data_log_force[7161] <= 16'h0000;
      coeffs_in_data_log_force[7162] <= 16'h0000;
      coeffs_in_data_log_force[7163] <= 16'h0000;
      coeffs_in_data_log_force[7164] <= 16'h0000;
      coeffs_in_data_log_force[7165] <= 16'h0000;
      coeffs_in_data_log_force[7166] <= 16'h0000;
      coeffs_in_data_log_force[7167] <= 16'h0000;
      coeffs_in_data_log_force[7168] <= 16'h0000;
      coeffs_in_data_log_force[7169] <= 16'h0000;
      coeffs_in_data_log_force[7170] <= 16'h0000;
      coeffs_in_data_log_force[7171] <= 16'h0000;
      coeffs_in_data_log_force[7172] <= 16'h0000;
      coeffs_in_data_log_force[7173] <= 16'h0000;
      coeffs_in_data_log_force[7174] <= 16'h0000;
      coeffs_in_data_log_force[7175] <= 16'h0000;
      coeffs_in_data_log_force[7176] <= 16'h0000;
      coeffs_in_data_log_force[7177] <= 16'h0000;
      coeffs_in_data_log_force[7178] <= 16'h0000;
      coeffs_in_data_log_force[7179] <= 16'h0000;
      coeffs_in_data_log_force[7180] <= 16'h0000;
      coeffs_in_data_log_force[7181] <= 16'h0000;
      coeffs_in_data_log_force[7182] <= 16'h0000;
      coeffs_in_data_log_force[7183] <= 16'h0000;
      coeffs_in_data_log_force[7184] <= 16'h0000;
      coeffs_in_data_log_force[7185] <= 16'h0000;
      coeffs_in_data_log_force[7186] <= 16'h0000;
      coeffs_in_data_log_force[7187] <= 16'h0000;
      coeffs_in_data_log_force[7188] <= 16'h0000;
      coeffs_in_data_log_force[7189] <= 16'h0000;
      coeffs_in_data_log_force[7190] <= 16'h0000;
      coeffs_in_data_log_force[7191] <= 16'h0000;
      coeffs_in_data_log_force[7192] <= 16'h0000;
      coeffs_in_data_log_force[7193] <= 16'h0000;
      coeffs_in_data_log_force[7194] <= 16'h0000;
      coeffs_in_data_log_force[7195] <= 16'h0000;
      coeffs_in_data_log_force[7196] <= 16'h0000;
      coeffs_in_data_log_force[7197] <= 16'h0000;
      coeffs_in_data_log_force[7198] <= 16'h0000;
      coeffs_in_data_log_force[7199] <= 16'h0000;
      coeffs_in_data_log_force[7200] <= 16'h0000;
      coeffs_in_data_log_force[7201] <= 16'h0000;
      coeffs_in_data_log_force[7202] <= 16'h0000;
      coeffs_in_data_log_force[7203] <= 16'h0000;
      coeffs_in_data_log_force[7204] <= 16'h0000;
      coeffs_in_data_log_force[7205] <= 16'h0000;
      coeffs_in_data_log_force[7206] <= 16'h0000;
      coeffs_in_data_log_force[7207] <= 16'h0000;
      coeffs_in_data_log_force[7208] <= 16'h0000;
      coeffs_in_data_log_force[7209] <= 16'h0000;
      coeffs_in_data_log_force[7210] <= 16'h0000;
      coeffs_in_data_log_force[7211] <= 16'h0000;
      coeffs_in_data_log_force[7212] <= 16'h0000;
      coeffs_in_data_log_force[7213] <= 16'h0000;
      coeffs_in_data_log_force[7214] <= 16'h0000;
      coeffs_in_data_log_force[7215] <= 16'h0000;
      coeffs_in_data_log_force[7216] <= 16'h0000;
      coeffs_in_data_log_force[7217] <= 16'h0000;
      coeffs_in_data_log_force[7218] <= 16'h0000;
      coeffs_in_data_log_force[7219] <= 16'h0000;
      coeffs_in_data_log_force[7220] <= 16'h0000;
      coeffs_in_data_log_force[7221] <= 16'h0000;
      coeffs_in_data_log_force[7222] <= 16'h0000;
      coeffs_in_data_log_force[7223] <= 16'h0000;
      coeffs_in_data_log_force[7224] <= 16'h0000;
      coeffs_in_data_log_force[7225] <= 16'h0000;
      coeffs_in_data_log_force[7226] <= 16'h0000;
      coeffs_in_data_log_force[7227] <= 16'h0000;
      coeffs_in_data_log_force[7228] <= 16'h0000;
      coeffs_in_data_log_force[7229] <= 16'h0000;
      coeffs_in_data_log_force[7230] <= 16'h0000;
      coeffs_in_data_log_force[7231] <= 16'h0000;
      coeffs_in_data_log_force[7232] <= 16'h0000;
      coeffs_in_data_log_force[7233] <= 16'h0000;
      coeffs_in_data_log_force[7234] <= 16'h0000;
      coeffs_in_data_log_force[7235] <= 16'h0000;
      coeffs_in_data_log_force[7236] <= 16'h0000;
      coeffs_in_data_log_force[7237] <= 16'h0000;
      coeffs_in_data_log_force[7238] <= 16'h0000;
      coeffs_in_data_log_force[7239] <= 16'h0000;
      coeffs_in_data_log_force[7240] <= 16'h0000;
      coeffs_in_data_log_force[7241] <= 16'h0000;
      coeffs_in_data_log_force[7242] <= 16'h0000;
      coeffs_in_data_log_force[7243] <= 16'h0000;
      coeffs_in_data_log_force[7244] <= 16'h0000;
      coeffs_in_data_log_force[7245] <= 16'h0000;
      coeffs_in_data_log_force[7246] <= 16'h0000;
      coeffs_in_data_log_force[7247] <= 16'h0000;
      coeffs_in_data_log_force[7248] <= 16'h0000;
      coeffs_in_data_log_force[7249] <= 16'h0000;
      coeffs_in_data_log_force[7250] <= 16'h0000;
      coeffs_in_data_log_force[7251] <= 16'h0000;
      coeffs_in_data_log_force[7252] <= 16'h0000;
      coeffs_in_data_log_force[7253] <= 16'h0000;
      coeffs_in_data_log_force[7254] <= 16'h0000;
      coeffs_in_data_log_force[7255] <= 16'h0000;
      coeffs_in_data_log_force[7256] <= 16'h0000;
      coeffs_in_data_log_force[7257] <= 16'h0000;
      coeffs_in_data_log_force[7258] <= 16'h0000;
      coeffs_in_data_log_force[7259] <= 16'h0000;
      coeffs_in_data_log_force[7260] <= 16'h0000;
      coeffs_in_data_log_force[7261] <= 16'h0000;
      coeffs_in_data_log_force[7262] <= 16'h0000;
      coeffs_in_data_log_force[7263] <= 16'h0000;
      coeffs_in_data_log_force[7264] <= 16'h0000;
      coeffs_in_data_log_force[7265] <= 16'h0000;
      coeffs_in_data_log_force[7266] <= 16'h0000;
      coeffs_in_data_log_force[7267] <= 16'h0000;
      coeffs_in_data_log_force[7268] <= 16'h0000;
      coeffs_in_data_log_force[7269] <= 16'h0000;
      coeffs_in_data_log_force[7270] <= 16'h0000;
      coeffs_in_data_log_force[7271] <= 16'h0000;
      coeffs_in_data_log_force[7272] <= 16'h0000;
      coeffs_in_data_log_force[7273] <= 16'h0000;
      coeffs_in_data_log_force[7274] <= 16'h0000;
      coeffs_in_data_log_force[7275] <= 16'h0000;
      coeffs_in_data_log_force[7276] <= 16'h0000;
      coeffs_in_data_log_force[7277] <= 16'h0000;
      coeffs_in_data_log_force[7278] <= 16'h0000;
      coeffs_in_data_log_force[7279] <= 16'h0000;
      coeffs_in_data_log_force[7280] <= 16'h0000;
      coeffs_in_data_log_force[7281] <= 16'h0000;
      coeffs_in_data_log_force[7282] <= 16'h0000;
      coeffs_in_data_log_force[7283] <= 16'h0000;
      coeffs_in_data_log_force[7284] <= 16'h0000;
      coeffs_in_data_log_force[7285] <= 16'h0000;
      coeffs_in_data_log_force[7286] <= 16'h0000;
      coeffs_in_data_log_force[7287] <= 16'h0000;
      coeffs_in_data_log_force[7288] <= 16'h0000;
      coeffs_in_data_log_force[7289] <= 16'h0000;
      coeffs_in_data_log_force[7290] <= 16'h0000;
      coeffs_in_data_log_force[7291] <= 16'h0000;
      coeffs_in_data_log_force[7292] <= 16'h0000;
      coeffs_in_data_log_force[7293] <= 16'h0000;
      coeffs_in_data_log_force[7294] <= 16'h0000;
      coeffs_in_data_log_force[7295] <= 16'h0000;
      coeffs_in_data_log_force[7296] <= 16'h0000;
      coeffs_in_data_log_force[7297] <= 16'h0000;
      coeffs_in_data_log_force[7298] <= 16'h0000;
      coeffs_in_data_log_force[7299] <= 16'h0000;
      coeffs_in_data_log_force[7300] <= 16'h0000;
      coeffs_in_data_log_force[7301] <= 16'h0000;
      coeffs_in_data_log_force[7302] <= 16'h0000;
      coeffs_in_data_log_force[7303] <= 16'h0000;
      coeffs_in_data_log_force[7304] <= 16'h0000;
      coeffs_in_data_log_force[7305] <= 16'h0000;
      coeffs_in_data_log_force[7306] <= 16'h0000;
      coeffs_in_data_log_force[7307] <= 16'h0000;
      coeffs_in_data_log_force[7308] <= 16'h0000;
      coeffs_in_data_log_force[7309] <= 16'h0000;
      coeffs_in_data_log_force[7310] <= 16'h0000;
      coeffs_in_data_log_force[7311] <= 16'h0000;
      coeffs_in_data_log_force[7312] <= 16'h0000;
      coeffs_in_data_log_force[7313] <= 16'h0000;
      coeffs_in_data_log_force[7314] <= 16'h0000;
      coeffs_in_data_log_force[7315] <= 16'h0000;
      coeffs_in_data_log_force[7316] <= 16'h0000;
      coeffs_in_data_log_force[7317] <= 16'h0000;
      coeffs_in_data_log_force[7318] <= 16'h0000;
      coeffs_in_data_log_force[7319] <= 16'h0000;
      coeffs_in_data_log_force[7320] <= 16'h0000;
      coeffs_in_data_log_force[7321] <= 16'h0000;
      coeffs_in_data_log_force[7322] <= 16'h0000;
      coeffs_in_data_log_force[7323] <= 16'h0000;
      coeffs_in_data_log_force[7324] <= 16'h0000;
      coeffs_in_data_log_force[7325] <= 16'h0000;
      coeffs_in_data_log_force[7326] <= 16'h0000;
      coeffs_in_data_log_force[7327] <= 16'h0000;
      coeffs_in_data_log_force[7328] <= 16'h0000;
      coeffs_in_data_log_force[7329] <= 16'h0000;
      coeffs_in_data_log_force[7330] <= 16'h0000;
      coeffs_in_data_log_force[7331] <= 16'h0000;
      coeffs_in_data_log_force[7332] <= 16'h0000;
      coeffs_in_data_log_force[7333] <= 16'h0000;
      coeffs_in_data_log_force[7334] <= 16'h0000;
      coeffs_in_data_log_force[7335] <= 16'h0000;
      coeffs_in_data_log_force[7336] <= 16'h0000;
      coeffs_in_data_log_force[7337] <= 16'h0000;
      coeffs_in_data_log_force[7338] <= 16'h0000;
      coeffs_in_data_log_force[7339] <= 16'h0000;
      coeffs_in_data_log_force[7340] <= 16'h0000;
      coeffs_in_data_log_force[7341] <= 16'h0000;
      coeffs_in_data_log_force[7342] <= 16'h0000;
      coeffs_in_data_log_force[7343] <= 16'h0000;
      coeffs_in_data_log_force[7344] <= 16'h0000;
      coeffs_in_data_log_force[7345] <= 16'h0000;
      coeffs_in_data_log_force[7346] <= 16'h0000;
      coeffs_in_data_log_force[7347] <= 16'h0000;
      coeffs_in_data_log_force[7348] <= 16'h0000;
      coeffs_in_data_log_force[7349] <= 16'h0000;
      coeffs_in_data_log_force[7350] <= 16'h0000;
      coeffs_in_data_log_force[7351] <= 16'h0000;
      coeffs_in_data_log_force[7352] <= 16'h0000;
      coeffs_in_data_log_force[7353] <= 16'h0000;
      coeffs_in_data_log_force[7354] <= 16'h0000;
      coeffs_in_data_log_force[7355] <= 16'h0000;
      coeffs_in_data_log_force[7356] <= 16'h0000;
      coeffs_in_data_log_force[7357] <= 16'h0000;
      coeffs_in_data_log_force[7358] <= 16'h0000;
      coeffs_in_data_log_force[7359] <= 16'h0000;
      coeffs_in_data_log_force[7360] <= 16'h0000;
      coeffs_in_data_log_force[7361] <= 16'h0000;
      coeffs_in_data_log_force[7362] <= 16'h0000;
      coeffs_in_data_log_force[7363] <= 16'h0000;
      coeffs_in_data_log_force[7364] <= 16'h0000;
      coeffs_in_data_log_force[7365] <= 16'h0000;
      coeffs_in_data_log_force[7366] <= 16'h0000;
      coeffs_in_data_log_force[7367] <= 16'h0000;
      coeffs_in_data_log_force[7368] <= 16'h0000;
      coeffs_in_data_log_force[7369] <= 16'h0000;
      coeffs_in_data_log_force[7370] <= 16'h0000;
      coeffs_in_data_log_force[7371] <= 16'h0000;
      coeffs_in_data_log_force[7372] <= 16'h0000;
      coeffs_in_data_log_force[7373] <= 16'h0000;
      coeffs_in_data_log_force[7374] <= 16'h0000;
      coeffs_in_data_log_force[7375] <= 16'h0000;
      coeffs_in_data_log_force[7376] <= 16'h0000;
      coeffs_in_data_log_force[7377] <= 16'h0000;
      coeffs_in_data_log_force[7378] <= 16'h0000;
      coeffs_in_data_log_force[7379] <= 16'h0000;
      coeffs_in_data_log_force[7380] <= 16'h0000;
      coeffs_in_data_log_force[7381] <= 16'h0000;
      coeffs_in_data_log_force[7382] <= 16'h0000;
      coeffs_in_data_log_force[7383] <= 16'h0000;
      coeffs_in_data_log_force[7384] <= 16'h0000;
      coeffs_in_data_log_force[7385] <= 16'h0000;
      coeffs_in_data_log_force[7386] <= 16'h0000;
      coeffs_in_data_log_force[7387] <= 16'h0000;
      coeffs_in_data_log_force[7388] <= 16'h0000;
      coeffs_in_data_log_force[7389] <= 16'h0000;
      coeffs_in_data_log_force[7390] <= 16'h0000;
      coeffs_in_data_log_force[7391] <= 16'h0000;
      coeffs_in_data_log_force[7392] <= 16'h0000;
      coeffs_in_data_log_force[7393] <= 16'h0000;
      coeffs_in_data_log_force[7394] <= 16'h0000;
      coeffs_in_data_log_force[7395] <= 16'h0000;
      coeffs_in_data_log_force[7396] <= 16'h0000;
      coeffs_in_data_log_force[7397] <= 16'h0000;
      coeffs_in_data_log_force[7398] <= 16'h0000;
      coeffs_in_data_log_force[7399] <= 16'h0000;
      coeffs_in_data_log_force[7400] <= 16'h0000;
      coeffs_in_data_log_force[7401] <= 16'h0000;
      coeffs_in_data_log_force[7402] <= 16'h0000;
      coeffs_in_data_log_force[7403] <= 16'h0000;
      coeffs_in_data_log_force[7404] <= 16'h0000;
      coeffs_in_data_log_force[7405] <= 16'h0000;
      coeffs_in_data_log_force[7406] <= 16'h0000;
      coeffs_in_data_log_force[7407] <= 16'h0000;
      coeffs_in_data_log_force[7408] <= 16'h0000;
      coeffs_in_data_log_force[7409] <= 16'h0000;
      coeffs_in_data_log_force[7410] <= 16'h0000;
      coeffs_in_data_log_force[7411] <= 16'h0000;
      coeffs_in_data_log_force[7412] <= 16'h0000;
      coeffs_in_data_log_force[7413] <= 16'h0000;
      coeffs_in_data_log_force[7414] <= 16'h0000;
      coeffs_in_data_log_force[7415] <= 16'h0000;
      coeffs_in_data_log_force[7416] <= 16'h0000;
      coeffs_in_data_log_force[7417] <= 16'h0000;
      coeffs_in_data_log_force[7418] <= 16'h0000;
      coeffs_in_data_log_force[7419] <= 16'h0000;
      coeffs_in_data_log_force[7420] <= 16'h0000;
      coeffs_in_data_log_force[7421] <= 16'h0000;
      coeffs_in_data_log_force[7422] <= 16'h0000;
      coeffs_in_data_log_force[7423] <= 16'h0000;
      coeffs_in_data_log_force[7424] <= 16'h0000;
      coeffs_in_data_log_force[7425] <= 16'h0000;
      coeffs_in_data_log_force[7426] <= 16'h0000;
      coeffs_in_data_log_force[7427] <= 16'h0000;
      coeffs_in_data_log_force[7428] <= 16'h0000;
      coeffs_in_data_log_force[7429] <= 16'h0000;
      coeffs_in_data_log_force[7430] <= 16'h0000;
      coeffs_in_data_log_force[7431] <= 16'h0000;
      coeffs_in_data_log_force[7432] <= 16'h0000;
      coeffs_in_data_log_force[7433] <= 16'h0000;
      coeffs_in_data_log_force[7434] <= 16'h0000;
      coeffs_in_data_log_force[7435] <= 16'h0000;
      coeffs_in_data_log_force[7436] <= 16'h0000;
      coeffs_in_data_log_force[7437] <= 16'h0000;
      coeffs_in_data_log_force[7438] <= 16'h0000;
      coeffs_in_data_log_force[7439] <= 16'h0000;
      coeffs_in_data_log_force[7440] <= 16'h0000;
      coeffs_in_data_log_force[7441] <= 16'h0000;
      coeffs_in_data_log_force[7442] <= 16'h0000;
      coeffs_in_data_log_force[7443] <= 16'h0000;
      coeffs_in_data_log_force[7444] <= 16'h0000;
      coeffs_in_data_log_force[7445] <= 16'h0000;
      coeffs_in_data_log_force[7446] <= 16'h0000;
      coeffs_in_data_log_force[7447] <= 16'h0000;
      coeffs_in_data_log_force[7448] <= 16'h0000;
      coeffs_in_data_log_force[7449] <= 16'h0000;
      coeffs_in_data_log_force[7450] <= 16'h0000;
      coeffs_in_data_log_force[7451] <= 16'h0000;
      coeffs_in_data_log_force[7452] <= 16'h0000;
      coeffs_in_data_log_force[7453] <= 16'h0000;
      coeffs_in_data_log_force[7454] <= 16'h0000;
      coeffs_in_data_log_force[7455] <= 16'h0000;
      coeffs_in_data_log_force[7456] <= 16'h0000;
      coeffs_in_data_log_force[7457] <= 16'h0000;
      coeffs_in_data_log_force[7458] <= 16'h0000;
      coeffs_in_data_log_force[7459] <= 16'h0000;
      coeffs_in_data_log_force[7460] <= 16'h0000;
      coeffs_in_data_log_force[7461] <= 16'h0000;
      coeffs_in_data_log_force[7462] <= 16'h0000;
      coeffs_in_data_log_force[7463] <= 16'h0000;
      coeffs_in_data_log_force[7464] <= 16'h0000;
      coeffs_in_data_log_force[7465] <= 16'h0000;
      coeffs_in_data_log_force[7466] <= 16'h0000;
      coeffs_in_data_log_force[7467] <= 16'h0000;
      coeffs_in_data_log_force[7468] <= 16'h0000;
      coeffs_in_data_log_force[7469] <= 16'h0000;
      coeffs_in_data_log_force[7470] <= 16'h0000;
      coeffs_in_data_log_force[7471] <= 16'h0000;
      coeffs_in_data_log_force[7472] <= 16'h0000;
      coeffs_in_data_log_force[7473] <= 16'h0000;
      coeffs_in_data_log_force[7474] <= 16'h0000;
      coeffs_in_data_log_force[7475] <= 16'h0000;
      coeffs_in_data_log_force[7476] <= 16'h0000;
      coeffs_in_data_log_force[7477] <= 16'h0000;
      coeffs_in_data_log_force[7478] <= 16'h0000;
      coeffs_in_data_log_force[7479] <= 16'h0000;
      coeffs_in_data_log_force[7480] <= 16'h0000;
      coeffs_in_data_log_force[7481] <= 16'h0000;
      coeffs_in_data_log_force[7482] <= 16'h0000;
      coeffs_in_data_log_force[7483] <= 16'h0000;
      coeffs_in_data_log_force[7484] <= 16'h0000;
      coeffs_in_data_log_force[7485] <= 16'h0000;
      coeffs_in_data_log_force[7486] <= 16'h0000;
      coeffs_in_data_log_force[7487] <= 16'h0000;
      coeffs_in_data_log_force[7488] <= 16'h0000;
      coeffs_in_data_log_force[7489] <= 16'h0000;
      coeffs_in_data_log_force[7490] <= 16'h0000;
      coeffs_in_data_log_force[7491] <= 16'h0000;
      coeffs_in_data_log_force[7492] <= 16'h0000;
      coeffs_in_data_log_force[7493] <= 16'h0000;
      coeffs_in_data_log_force[7494] <= 16'h0000;
      coeffs_in_data_log_force[7495] <= 16'h0000;
      coeffs_in_data_log_force[7496] <= 16'h0000;
      coeffs_in_data_log_force[7497] <= 16'h0000;
      coeffs_in_data_log_force[7498] <= 16'h0000;
      coeffs_in_data_log_force[7499] <= 16'h0000;
      coeffs_in_data_log_force[7500] <= 16'h0000;
      coeffs_in_data_log_force[7501] <= 16'h0000;
      coeffs_in_data_log_force[7502] <= 16'h0000;
      coeffs_in_data_log_force[7503] <= 16'h0000;
      coeffs_in_data_log_force[7504] <= 16'h0000;
      coeffs_in_data_log_force[7505] <= 16'h0000;
      coeffs_in_data_log_force[7506] <= 16'h0000;
      coeffs_in_data_log_force[7507] <= 16'h0000;
      coeffs_in_data_log_force[7508] <= 16'h0000;
      coeffs_in_data_log_force[7509] <= 16'h0000;
      coeffs_in_data_log_force[7510] <= 16'h0000;
      coeffs_in_data_log_force[7511] <= 16'h0000;
      coeffs_in_data_log_force[7512] <= 16'h0000;
      coeffs_in_data_log_force[7513] <= 16'h0000;
      coeffs_in_data_log_force[7514] <= 16'h0000;
      coeffs_in_data_log_force[7515] <= 16'h0000;
      coeffs_in_data_log_force[7516] <= 16'h0000;
      coeffs_in_data_log_force[7517] <= 16'h0000;
      coeffs_in_data_log_force[7518] <= 16'h0000;
      coeffs_in_data_log_force[7519] <= 16'h0000;
      coeffs_in_data_log_force[7520] <= 16'h0000;
      coeffs_in_data_log_force[7521] <= 16'h0000;
      coeffs_in_data_log_force[7522] <= 16'h0000;
      coeffs_in_data_log_force[7523] <= 16'h0000;
      coeffs_in_data_log_force[7524] <= 16'h0000;
      coeffs_in_data_log_force[7525] <= 16'h0000;
      coeffs_in_data_log_force[7526] <= 16'h0000;
      coeffs_in_data_log_force[7527] <= 16'h0000;
      coeffs_in_data_log_force[7528] <= 16'h0000;
      coeffs_in_data_log_force[7529] <= 16'h0000;
      coeffs_in_data_log_force[7530] <= 16'h0000;
      coeffs_in_data_log_force[7531] <= 16'h0000;
      coeffs_in_data_log_force[7532] <= 16'h0000;
      coeffs_in_data_log_force[7533] <= 16'h0000;
      coeffs_in_data_log_force[7534] <= 16'h0000;
      coeffs_in_data_log_force[7535] <= 16'h0000;
      coeffs_in_data_log_force[7536] <= 16'h0000;
      coeffs_in_data_log_force[7537] <= 16'h0000;
      coeffs_in_data_log_force[7538] <= 16'h0000;
      coeffs_in_data_log_force[7539] <= 16'h0000;
      coeffs_in_data_log_force[7540] <= 16'h0000;
      coeffs_in_data_log_force[7541] <= 16'h0000;
      coeffs_in_data_log_force[7542] <= 16'h0000;
      coeffs_in_data_log_force[7543] <= 16'h0000;
      coeffs_in_data_log_force[7544] <= 16'h0000;
      coeffs_in_data_log_force[7545] <= 16'h0000;
      coeffs_in_data_log_force[7546] <= 16'h0000;
      coeffs_in_data_log_force[7547] <= 16'h0000;
      coeffs_in_data_log_force[7548] <= 16'h0000;
      coeffs_in_data_log_force[7549] <= 16'h0000;
      coeffs_in_data_log_force[7550] <= 16'h0000;
      coeffs_in_data_log_force[7551] <= 16'h0000;
      coeffs_in_data_log_force[7552] <= 16'h0000;
      coeffs_in_data_log_force[7553] <= 16'h0000;
      coeffs_in_data_log_force[7554] <= 16'h0000;
      coeffs_in_data_log_force[7555] <= 16'h0000;
      coeffs_in_data_log_force[7556] <= 16'h0000;
      coeffs_in_data_log_force[7557] <= 16'h0000;
      coeffs_in_data_log_force[7558] <= 16'h0000;
      coeffs_in_data_log_force[7559] <= 16'h0000;
      coeffs_in_data_log_force[7560] <= 16'h0000;
      coeffs_in_data_log_force[7561] <= 16'h0000;
      coeffs_in_data_log_force[7562] <= 16'h0000;
      coeffs_in_data_log_force[7563] <= 16'h0000;
      coeffs_in_data_log_force[7564] <= 16'h0000;
      coeffs_in_data_log_force[7565] <= 16'h0000;
      coeffs_in_data_log_force[7566] <= 16'h0000;
      coeffs_in_data_log_force[7567] <= 16'h0000;
      coeffs_in_data_log_force[7568] <= 16'h0000;
      coeffs_in_data_log_force[7569] <= 16'h0000;
      coeffs_in_data_log_force[7570] <= 16'h0000;
      coeffs_in_data_log_force[7571] <= 16'h0000;
      coeffs_in_data_log_force[7572] <= 16'h0000;
      coeffs_in_data_log_force[7573] <= 16'h0000;
      coeffs_in_data_log_force[7574] <= 16'h0000;
      coeffs_in_data_log_force[7575] <= 16'h0000;
      coeffs_in_data_log_force[7576] <= 16'h0000;
      coeffs_in_data_log_force[7577] <= 16'h0000;
      coeffs_in_data_log_force[7578] <= 16'h0000;
      coeffs_in_data_log_force[7579] <= 16'h0000;
      coeffs_in_data_log_force[7580] <= 16'h0000;
      coeffs_in_data_log_force[7581] <= 16'h0000;
      coeffs_in_data_log_force[7582] <= 16'h0000;
      coeffs_in_data_log_force[7583] <= 16'h0000;
      coeffs_in_data_log_force[7584] <= 16'h0000;
      coeffs_in_data_log_force[7585] <= 16'h0000;
      coeffs_in_data_log_force[7586] <= 16'h0000;
      coeffs_in_data_log_force[7587] <= 16'h0000;
      coeffs_in_data_log_force[7588] <= 16'h0000;
      coeffs_in_data_log_force[7589] <= 16'h0000;
      coeffs_in_data_log_force[7590] <= 16'h0000;
      coeffs_in_data_log_force[7591] <= 16'h0000;
      coeffs_in_data_log_force[7592] <= 16'h0000;
      coeffs_in_data_log_force[7593] <= 16'h0000;
      coeffs_in_data_log_force[7594] <= 16'h0000;
      coeffs_in_data_log_force[7595] <= 16'h0000;
      coeffs_in_data_log_force[7596] <= 16'h0000;
      coeffs_in_data_log_force[7597] <= 16'h0000;
      coeffs_in_data_log_force[7598] <= 16'h0000;
      coeffs_in_data_log_force[7599] <= 16'h0000;
      coeffs_in_data_log_force[7600] <= 16'h0000;
      coeffs_in_data_log_force[7601] <= 16'h0000;
      coeffs_in_data_log_force[7602] <= 16'h0000;
      coeffs_in_data_log_force[7603] <= 16'h0000;
      coeffs_in_data_log_force[7604] <= 16'h0000;
      coeffs_in_data_log_force[7605] <= 16'h0000;
      coeffs_in_data_log_force[7606] <= 16'h0000;
      coeffs_in_data_log_force[7607] <= 16'h0000;
      coeffs_in_data_log_force[7608] <= 16'h0000;
      coeffs_in_data_log_force[7609] <= 16'h0000;
      coeffs_in_data_log_force[7610] <= 16'h0000;
      coeffs_in_data_log_force[7611] <= 16'h0000;
      coeffs_in_data_log_force[7612] <= 16'h0000;
      coeffs_in_data_log_force[7613] <= 16'h0000;
      coeffs_in_data_log_force[7614] <= 16'h0000;
      coeffs_in_data_log_force[7615] <= 16'h0000;
      coeffs_in_data_log_force[7616] <= 16'h0000;
      coeffs_in_data_log_force[7617] <= 16'h0000;
      coeffs_in_data_log_force[7618] <= 16'h0000;
      coeffs_in_data_log_force[7619] <= 16'h0000;
      coeffs_in_data_log_force[7620] <= 16'h0000;
      coeffs_in_data_log_force[7621] <= 16'h0000;
      coeffs_in_data_log_force[7622] <= 16'h0000;
      coeffs_in_data_log_force[7623] <= 16'h0000;
      coeffs_in_data_log_force[7624] <= 16'h0000;
      coeffs_in_data_log_force[7625] <= 16'h0000;
      coeffs_in_data_log_force[7626] <= 16'h0000;
      coeffs_in_data_log_force[7627] <= 16'h0000;
      coeffs_in_data_log_force[7628] <= 16'h0000;
      coeffs_in_data_log_force[7629] <= 16'h0000;
      coeffs_in_data_log_force[7630] <= 16'h0000;
      coeffs_in_data_log_force[7631] <= 16'h0000;
      coeffs_in_data_log_force[7632] <= 16'h0000;
      coeffs_in_data_log_force[7633] <= 16'h0000;
      coeffs_in_data_log_force[7634] <= 16'h0000;
      coeffs_in_data_log_force[7635] <= 16'h0000;
      coeffs_in_data_log_force[7636] <= 16'h0000;
      coeffs_in_data_log_force[7637] <= 16'h0000;
      coeffs_in_data_log_force[7638] <= 16'h0000;
      coeffs_in_data_log_force[7639] <= 16'h0000;
      coeffs_in_data_log_force[7640] <= 16'h0000;
      coeffs_in_data_log_force[7641] <= 16'h0000;
      coeffs_in_data_log_force[7642] <= 16'h0000;
      coeffs_in_data_log_force[7643] <= 16'h0000;
      coeffs_in_data_log_force[7644] <= 16'h0000;
      coeffs_in_data_log_force[7645] <= 16'h0000;
      coeffs_in_data_log_force[7646] <= 16'h0000;
      coeffs_in_data_log_force[7647] <= 16'h0000;
      coeffs_in_data_log_force[7648] <= 16'h0000;
      coeffs_in_data_log_force[7649] <= 16'h0000;
      coeffs_in_data_log_force[7650] <= 16'h0000;
      coeffs_in_data_log_force[7651] <= 16'h0000;
      coeffs_in_data_log_force[7652] <= 16'h0000;
      coeffs_in_data_log_force[7653] <= 16'h0000;
      coeffs_in_data_log_force[7654] <= 16'h0000;
      coeffs_in_data_log_force[7655] <= 16'h0000;
      coeffs_in_data_log_force[7656] <= 16'h0000;
      coeffs_in_data_log_force[7657] <= 16'h0000;
      coeffs_in_data_log_force[7658] <= 16'h0000;
      coeffs_in_data_log_force[7659] <= 16'h0000;
      coeffs_in_data_log_force[7660] <= 16'h0000;
      coeffs_in_data_log_force[7661] <= 16'h0000;
      coeffs_in_data_log_force[7662] <= 16'h0000;
      coeffs_in_data_log_force[7663] <= 16'h0000;
      coeffs_in_data_log_force[7664] <= 16'h0000;
      coeffs_in_data_log_force[7665] <= 16'h0000;
      coeffs_in_data_log_force[7666] <= 16'h0000;
      coeffs_in_data_log_force[7667] <= 16'h0000;
      coeffs_in_data_log_force[7668] <= 16'h0000;
      coeffs_in_data_log_force[7669] <= 16'h0000;
      coeffs_in_data_log_force[7670] <= 16'h0000;
      coeffs_in_data_log_force[7671] <= 16'h0000;
      coeffs_in_data_log_force[7672] <= 16'h0000;
      coeffs_in_data_log_force[7673] <= 16'h0000;
      coeffs_in_data_log_force[7674] <= 16'h0000;
      coeffs_in_data_log_force[7675] <= 16'h0000;
      coeffs_in_data_log_force[7676] <= 16'h0000;
      coeffs_in_data_log_force[7677] <= 16'h0000;
      coeffs_in_data_log_force[7678] <= 16'h0000;
      coeffs_in_data_log_force[7679] <= 16'h0000;
      coeffs_in_data_log_force[7680] <= 16'h0000;
      coeffs_in_data_log_force[7681] <= 16'h0000;
      coeffs_in_data_log_force[7682] <= 16'h0000;
      coeffs_in_data_log_force[7683] <= 16'h0000;
      coeffs_in_data_log_force[7684] <= 16'h0000;
      coeffs_in_data_log_force[7685] <= 16'h0000;
      coeffs_in_data_log_force[7686] <= 16'h0000;
      coeffs_in_data_log_force[7687] <= 16'h0000;
      coeffs_in_data_log_force[7688] <= 16'h0000;
      coeffs_in_data_log_force[7689] <= 16'h0000;
      coeffs_in_data_log_force[7690] <= 16'h0000;
      coeffs_in_data_log_force[7691] <= 16'h0000;
      coeffs_in_data_log_force[7692] <= 16'h0000;
      coeffs_in_data_log_force[7693] <= 16'h0000;
      coeffs_in_data_log_force[7694] <= 16'h0000;
      coeffs_in_data_log_force[7695] <= 16'h0000;
      coeffs_in_data_log_force[7696] <= 16'h0000;
      coeffs_in_data_log_force[7697] <= 16'h0000;
      coeffs_in_data_log_force[7698] <= 16'h0000;
      coeffs_in_data_log_force[7699] <= 16'h0000;
      coeffs_in_data_log_force[7700] <= 16'h0000;
      coeffs_in_data_log_force[7701] <= 16'h0000;
      coeffs_in_data_log_force[7702] <= 16'h0000;
      coeffs_in_data_log_force[7703] <= 16'h0000;
      coeffs_in_data_log_force[7704] <= 16'h0000;
      coeffs_in_data_log_force[7705] <= 16'h0000;
      coeffs_in_data_log_force[7706] <= 16'h0000;
      coeffs_in_data_log_force[7707] <= 16'h0000;
      coeffs_in_data_log_force[7708] <= 16'h0000;
      coeffs_in_data_log_force[7709] <= 16'h0000;
      coeffs_in_data_log_force[7710] <= 16'h0000;
      coeffs_in_data_log_force[7711] <= 16'h0000;
      coeffs_in_data_log_force[7712] <= 16'h0000;
      coeffs_in_data_log_force[7713] <= 16'h0000;
      coeffs_in_data_log_force[7714] <= 16'h0000;
      coeffs_in_data_log_force[7715] <= 16'h0000;
      coeffs_in_data_log_force[7716] <= 16'h0000;
      coeffs_in_data_log_force[7717] <= 16'h0000;
      coeffs_in_data_log_force[7718] <= 16'h0000;
      coeffs_in_data_log_force[7719] <= 16'h0000;
      coeffs_in_data_log_force[7720] <= 16'h0000;
      coeffs_in_data_log_force[7721] <= 16'h0000;
      coeffs_in_data_log_force[7722] <= 16'h0000;
      coeffs_in_data_log_force[7723] <= 16'h0000;
      coeffs_in_data_log_force[7724] <= 16'h0000;
      coeffs_in_data_log_force[7725] <= 16'h0000;
      coeffs_in_data_log_force[7726] <= 16'h0000;
      coeffs_in_data_log_force[7727] <= 16'h0000;
      coeffs_in_data_log_force[7728] <= 16'h0000;
      coeffs_in_data_log_force[7729] <= 16'h0000;
      coeffs_in_data_log_force[7730] <= 16'h0000;
      coeffs_in_data_log_force[7731] <= 16'h0000;
      coeffs_in_data_log_force[7732] <= 16'h0000;
      coeffs_in_data_log_force[7733] <= 16'h0000;
      coeffs_in_data_log_force[7734] <= 16'h0000;
      coeffs_in_data_log_force[7735] <= 16'h0000;
      coeffs_in_data_log_force[7736] <= 16'h0000;
      coeffs_in_data_log_force[7737] <= 16'h0000;
      coeffs_in_data_log_force[7738] <= 16'h0000;
      coeffs_in_data_log_force[7739] <= 16'h0000;
      coeffs_in_data_log_force[7740] <= 16'h0000;
      coeffs_in_data_log_force[7741] <= 16'h0000;
      coeffs_in_data_log_force[7742] <= 16'h0000;
      coeffs_in_data_log_force[7743] <= 16'h0000;
      coeffs_in_data_log_force[7744] <= 16'h0000;
      coeffs_in_data_log_force[7745] <= 16'h0000;
      coeffs_in_data_log_force[7746] <= 16'h0000;
      coeffs_in_data_log_force[7747] <= 16'h0000;
      coeffs_in_data_log_force[7748] <= 16'h0000;
      coeffs_in_data_log_force[7749] <= 16'h0000;
      coeffs_in_data_log_force[7750] <= 16'h0000;
      coeffs_in_data_log_force[7751] <= 16'h0000;
      coeffs_in_data_log_force[7752] <= 16'h0000;
      coeffs_in_data_log_force[7753] <= 16'h0000;
      coeffs_in_data_log_force[7754] <= 16'h0000;
      coeffs_in_data_log_force[7755] <= 16'h0000;
      coeffs_in_data_log_force[7756] <= 16'h0000;
      coeffs_in_data_log_force[7757] <= 16'h0000;
      coeffs_in_data_log_force[7758] <= 16'h0000;
      coeffs_in_data_log_force[7759] <= 16'h0000;
      coeffs_in_data_log_force[7760] <= 16'h0000;
      coeffs_in_data_log_force[7761] <= 16'h0000;
      coeffs_in_data_log_force[7762] <= 16'h0000;
      coeffs_in_data_log_force[7763] <= 16'h0000;
      coeffs_in_data_log_force[7764] <= 16'h0000;
      coeffs_in_data_log_force[7765] <= 16'h0000;
      coeffs_in_data_log_force[7766] <= 16'h0000;
      coeffs_in_data_log_force[7767] <= 16'h0000;
      coeffs_in_data_log_force[7768] <= 16'h0000;
      coeffs_in_data_log_force[7769] <= 16'h0000;
      coeffs_in_data_log_force[7770] <= 16'h0000;
      coeffs_in_data_log_force[7771] <= 16'h0000;
      coeffs_in_data_log_force[7772] <= 16'h0000;
      coeffs_in_data_log_force[7773] <= 16'h0000;
      coeffs_in_data_log_force[7774] <= 16'h0000;
      coeffs_in_data_log_force[7775] <= 16'h0000;
      coeffs_in_data_log_force[7776] <= 16'h0000;
      coeffs_in_data_log_force[7777] <= 16'h0000;
      coeffs_in_data_log_force[7778] <= 16'h0000;
      coeffs_in_data_log_force[7779] <= 16'h0000;
      coeffs_in_data_log_force[7780] <= 16'h0000;
      coeffs_in_data_log_force[7781] <= 16'h0000;
      coeffs_in_data_log_force[7782] <= 16'h0000;
      coeffs_in_data_log_force[7783] <= 16'h0000;
      coeffs_in_data_log_force[7784] <= 16'h0000;
      coeffs_in_data_log_force[7785] <= 16'h0000;
      coeffs_in_data_log_force[7786] <= 16'h0000;
      coeffs_in_data_log_force[7787] <= 16'h0000;
      coeffs_in_data_log_force[7788] <= 16'h0000;
      coeffs_in_data_log_force[7789] <= 16'h0000;
      coeffs_in_data_log_force[7790] <= 16'h0000;
      coeffs_in_data_log_force[7791] <= 16'h0000;
      coeffs_in_data_log_force[7792] <= 16'h0000;
      coeffs_in_data_log_force[7793] <= 16'h0000;
      coeffs_in_data_log_force[7794] <= 16'h0000;
      coeffs_in_data_log_force[7795] <= 16'h0000;
      coeffs_in_data_log_force[7796] <= 16'h0000;
      coeffs_in_data_log_force[7797] <= 16'h0000;
      coeffs_in_data_log_force[7798] <= 16'h0000;
      coeffs_in_data_log_force[7799] <= 16'h0000;
      coeffs_in_data_log_force[7800] <= 16'h0000;
      coeffs_in_data_log_force[7801] <= 16'h0000;
      coeffs_in_data_log_force[7802] <= 16'h0000;
      coeffs_in_data_log_force[7803] <= 16'h0000;
      coeffs_in_data_log_force[7804] <= 16'h0000;
      coeffs_in_data_log_force[7805] <= 16'h0000;
      coeffs_in_data_log_force[7806] <= 16'h0000;
      coeffs_in_data_log_force[7807] <= 16'h0000;
      coeffs_in_data_log_force[7808] <= 16'h0000;
      coeffs_in_data_log_force[7809] <= 16'h0000;
      coeffs_in_data_log_force[7810] <= 16'h0000;
      coeffs_in_data_log_force[7811] <= 16'h0000;
      coeffs_in_data_log_force[7812] <= 16'h0000;
      coeffs_in_data_log_force[7813] <= 16'h0000;
      coeffs_in_data_log_force[7814] <= 16'h0000;
      coeffs_in_data_log_force[7815] <= 16'h0000;
      coeffs_in_data_log_force[7816] <= 16'h0000;
      coeffs_in_data_log_force[7817] <= 16'h0000;
      coeffs_in_data_log_force[7818] <= 16'h0000;
      coeffs_in_data_log_force[7819] <= 16'h0000;
      coeffs_in_data_log_force[7820] <= 16'h0000;
      coeffs_in_data_log_force[7821] <= 16'h0000;
      coeffs_in_data_log_force[7822] <= 16'h0000;
      coeffs_in_data_log_force[7823] <= 16'h0000;
      coeffs_in_data_log_force[7824] <= 16'h0000;
      coeffs_in_data_log_force[7825] <= 16'h0000;
      coeffs_in_data_log_force[7826] <= 16'h0000;
      coeffs_in_data_log_force[7827] <= 16'h0000;
      coeffs_in_data_log_force[7828] <= 16'h0000;
      coeffs_in_data_log_force[7829] <= 16'h0000;
      coeffs_in_data_log_force[7830] <= 16'h0000;
      coeffs_in_data_log_force[7831] <= 16'h0000;
      coeffs_in_data_log_force[7832] <= 16'h0000;
      coeffs_in_data_log_force[7833] <= 16'h0000;
      coeffs_in_data_log_force[7834] <= 16'h0000;
      coeffs_in_data_log_force[7835] <= 16'h0000;
      coeffs_in_data_log_force[7836] <= 16'h0000;
      coeffs_in_data_log_force[7837] <= 16'h0000;
      coeffs_in_data_log_force[7838] <= 16'h0000;
      coeffs_in_data_log_force[7839] <= 16'h0000;
      coeffs_in_data_log_force[7840] <= 16'h0000;
      coeffs_in_data_log_force[7841] <= 16'h0000;
      coeffs_in_data_log_force[7842] <= 16'h0000;
      coeffs_in_data_log_force[7843] <= 16'h0000;
      coeffs_in_data_log_force[7844] <= 16'h0000;
      coeffs_in_data_log_force[7845] <= 16'h0000;
      coeffs_in_data_log_force[7846] <= 16'h0000;
      coeffs_in_data_log_force[7847] <= 16'h0000;
      coeffs_in_data_log_force[7848] <= 16'h0000;
      coeffs_in_data_log_force[7849] <= 16'h0000;
      coeffs_in_data_log_force[7850] <= 16'h0000;
      coeffs_in_data_log_force[7851] <= 16'h0000;
      coeffs_in_data_log_force[7852] <= 16'h0000;
      coeffs_in_data_log_force[7853] <= 16'h0000;
      coeffs_in_data_log_force[7854] <= 16'h0000;
      coeffs_in_data_log_force[7855] <= 16'h0000;
      coeffs_in_data_log_force[7856] <= 16'h0000;
      coeffs_in_data_log_force[7857] <= 16'h0000;
      coeffs_in_data_log_force[7858] <= 16'h0000;
      coeffs_in_data_log_force[7859] <= 16'h0000;
      coeffs_in_data_log_force[7860] <= 16'h0000;
      coeffs_in_data_log_force[7861] <= 16'h0000;
      coeffs_in_data_log_force[7862] <= 16'h0000;
      coeffs_in_data_log_force[7863] <= 16'h0000;
      coeffs_in_data_log_force[7864] <= 16'h0000;
      coeffs_in_data_log_force[7865] <= 16'h0000;
      coeffs_in_data_log_force[7866] <= 16'h0000;
      coeffs_in_data_log_force[7867] <= 16'h0000;
      coeffs_in_data_log_force[7868] <= 16'h0000;
      coeffs_in_data_log_force[7869] <= 16'h0000;
      coeffs_in_data_log_force[7870] <= 16'h0000;
      coeffs_in_data_log_force[7871] <= 16'h0000;
      coeffs_in_data_log_force[7872] <= 16'h0000;
      coeffs_in_data_log_force[7873] <= 16'h0000;
      coeffs_in_data_log_force[7874] <= 16'h0000;
      coeffs_in_data_log_force[7875] <= 16'h0000;
      coeffs_in_data_log_force[7876] <= 16'h0000;
      coeffs_in_data_log_force[7877] <= 16'h0000;
      coeffs_in_data_log_force[7878] <= 16'h0000;
      coeffs_in_data_log_force[7879] <= 16'h0000;
      coeffs_in_data_log_force[7880] <= 16'h0000;
      coeffs_in_data_log_force[7881] <= 16'h0000;
      coeffs_in_data_log_force[7882] <= 16'h0000;
      coeffs_in_data_log_force[7883] <= 16'h0000;
      coeffs_in_data_log_force[7884] <= 16'h0000;
      coeffs_in_data_log_force[7885] <= 16'h0000;
      coeffs_in_data_log_force[7886] <= 16'h0000;
      coeffs_in_data_log_force[7887] <= 16'h0000;
      coeffs_in_data_log_force[7888] <= 16'h0000;
      coeffs_in_data_log_force[7889] <= 16'h0000;
      coeffs_in_data_log_force[7890] <= 16'h0000;
      coeffs_in_data_log_force[7891] <= 16'h0000;
      coeffs_in_data_log_force[7892] <= 16'h0000;
      coeffs_in_data_log_force[7893] <= 16'h0000;
      coeffs_in_data_log_force[7894] <= 16'h0000;
      coeffs_in_data_log_force[7895] <= 16'h0000;
      coeffs_in_data_log_force[7896] <= 16'h0000;
      coeffs_in_data_log_force[7897] <= 16'h0000;
      coeffs_in_data_log_force[7898] <= 16'h0000;
      coeffs_in_data_log_force[7899] <= 16'h0000;
      coeffs_in_data_log_force[7900] <= 16'h0000;
      coeffs_in_data_log_force[7901] <= 16'h0000;
      coeffs_in_data_log_force[7902] <= 16'h0000;
      coeffs_in_data_log_force[7903] <= 16'h0000;
      coeffs_in_data_log_force[7904] <= 16'h0000;
      coeffs_in_data_log_force[7905] <= 16'h0000;
      coeffs_in_data_log_force[7906] <= 16'h0000;
      coeffs_in_data_log_force[7907] <= 16'h0000;
      coeffs_in_data_log_force[7908] <= 16'h0000;
      coeffs_in_data_log_force[7909] <= 16'h0000;
      coeffs_in_data_log_force[7910] <= 16'h0000;
      coeffs_in_data_log_force[7911] <= 16'h0000;
      coeffs_in_data_log_force[7912] <= 16'h0000;
      coeffs_in_data_log_force[7913] <= 16'h0000;
      coeffs_in_data_log_force[7914] <= 16'h0000;
      coeffs_in_data_log_force[7915] <= 16'h0000;
      coeffs_in_data_log_force[7916] <= 16'h0000;
      coeffs_in_data_log_force[7917] <= 16'h0000;
      coeffs_in_data_log_force[7918] <= 16'h0000;
      coeffs_in_data_log_force[7919] <= 16'h0000;
      coeffs_in_data_log_force[7920] <= 16'h0000;
      coeffs_in_data_log_force[7921] <= 16'h0000;
      coeffs_in_data_log_force[7922] <= 16'h0000;
      coeffs_in_data_log_force[7923] <= 16'h0000;
      coeffs_in_data_log_force[7924] <= 16'h0000;
      coeffs_in_data_log_force[7925] <= 16'h0000;
      coeffs_in_data_log_force[7926] <= 16'h0000;
      coeffs_in_data_log_force[7927] <= 16'h0000;
      coeffs_in_data_log_force[7928] <= 16'h0000;
      coeffs_in_data_log_force[7929] <= 16'h0000;
      coeffs_in_data_log_force[7930] <= 16'h0000;
      coeffs_in_data_log_force[7931] <= 16'h0000;
      coeffs_in_data_log_force[7932] <= 16'h0000;
      coeffs_in_data_log_force[7933] <= 16'h0000;
      coeffs_in_data_log_force[7934] <= 16'h0000;
      coeffs_in_data_log_force[7935] <= 16'h0000;
      coeffs_in_data_log_force[7936] <= 16'h0000;
      coeffs_in_data_log_force[7937] <= 16'h0000;
      coeffs_in_data_log_force[7938] <= 16'h0000;
      coeffs_in_data_log_force[7939] <= 16'h0000;
      coeffs_in_data_log_force[7940] <= 16'h0000;
      coeffs_in_data_log_force[7941] <= 16'h0000;
      coeffs_in_data_log_force[7942] <= 16'h0000;
      coeffs_in_data_log_force[7943] <= 16'h0000;
      coeffs_in_data_log_force[7944] <= 16'h0000;
      coeffs_in_data_log_force[7945] <= 16'h0000;
      coeffs_in_data_log_force[7946] <= 16'h0000;
      coeffs_in_data_log_force[7947] <= 16'h0000;
      coeffs_in_data_log_force[7948] <= 16'h0000;
      coeffs_in_data_log_force[7949] <= 16'h0000;
      coeffs_in_data_log_force[7950] <= 16'h0000;
      coeffs_in_data_log_force[7951] <= 16'h0000;
      coeffs_in_data_log_force[7952] <= 16'h0000;
      coeffs_in_data_log_force[7953] <= 16'h0000;
      coeffs_in_data_log_force[7954] <= 16'h0000;
      coeffs_in_data_log_force[7955] <= 16'h0000;
      coeffs_in_data_log_force[7956] <= 16'h0000;
      coeffs_in_data_log_force[7957] <= 16'h0000;
      coeffs_in_data_log_force[7958] <= 16'h0000;
      coeffs_in_data_log_force[7959] <= 16'h0000;
      coeffs_in_data_log_force[7960] <= 16'h0000;
      coeffs_in_data_log_force[7961] <= 16'h0000;
      coeffs_in_data_log_force[7962] <= 16'h0000;
      coeffs_in_data_log_force[7963] <= 16'h0000;
      coeffs_in_data_log_force[7964] <= 16'h0000;
      coeffs_in_data_log_force[7965] <= 16'h0000;
      coeffs_in_data_log_force[7966] <= 16'h0000;
      coeffs_in_data_log_force[7967] <= 16'h0000;
      coeffs_in_data_log_force[7968] <= 16'h0000;
      coeffs_in_data_log_force[7969] <= 16'h0000;
      coeffs_in_data_log_force[7970] <= 16'h0000;
      coeffs_in_data_log_force[7971] <= 16'h0000;
      coeffs_in_data_log_force[7972] <= 16'h0000;
      coeffs_in_data_log_force[7973] <= 16'h0000;
      coeffs_in_data_log_force[7974] <= 16'h0000;
      coeffs_in_data_log_force[7975] <= 16'h0000;
      coeffs_in_data_log_force[7976] <= 16'h0000;
      coeffs_in_data_log_force[7977] <= 16'h0000;
      coeffs_in_data_log_force[7978] <= 16'h0000;
      coeffs_in_data_log_force[7979] <= 16'h0000;
      coeffs_in_data_log_force[7980] <= 16'h0000;
      coeffs_in_data_log_force[7981] <= 16'h0000;
      coeffs_in_data_log_force[7982] <= 16'h0000;
      coeffs_in_data_log_force[7983] <= 16'h0000;
      coeffs_in_data_log_force[7984] <= 16'h0000;
      coeffs_in_data_log_force[7985] <= 16'h0000;
      coeffs_in_data_log_force[7986] <= 16'h0000;
      coeffs_in_data_log_force[7987] <= 16'h0000;
      coeffs_in_data_log_force[7988] <= 16'h0000;
      coeffs_in_data_log_force[7989] <= 16'h0000;
      coeffs_in_data_log_force[7990] <= 16'h0000;
      coeffs_in_data_log_force[7991] <= 16'h0000;
      coeffs_in_data_log_force[7992] <= 16'h0000;
      coeffs_in_data_log_force[7993] <= 16'h0000;
      coeffs_in_data_log_force[7994] <= 16'h0000;
      coeffs_in_data_log_force[7995] <= 16'h0000;
      coeffs_in_data_log_force[7996] <= 16'h0000;
      coeffs_in_data_log_force[7997] <= 16'h0000;
      coeffs_in_data_log_force[7998] <= 16'h0000;
      coeffs_in_data_log_force[7999] <= 16'h0000;
      coeffs_in_data_log_force[8000] <= 16'h0000;
      coeffs_in_data_log_force[8001] <= 16'h0000;
      coeffs_in_data_log_force[8002] <= 16'h0000;
      coeffs_in_data_log_force[8003] <= 16'h0000;
      coeffs_in_data_log_force[8004] <= 16'h0000;
      coeffs_in_data_log_force[8005] <= 16'h0000;
      coeffs_in_data_log_force[8006] <= 16'h0000;
      coeffs_in_data_log_force[8007] <= 16'h0000;
      coeffs_in_data_log_force[8008] <= 16'h0000;
      coeffs_in_data_log_force[8009] <= 16'h0000;
      coeffs_in_data_log_force[8010] <= 16'h0000;
      coeffs_in_data_log_force[8011] <= 16'h0000;
      coeffs_in_data_log_force[8012] <= 16'h0000;
      coeffs_in_data_log_force[8013] <= 16'h0000;
      coeffs_in_data_log_force[8014] <= 16'h0000;
      coeffs_in_data_log_force[8015] <= 16'h0000;
      coeffs_in_data_log_force[8016] <= 16'h0000;
      coeffs_in_data_log_force[8017] <= 16'h0000;
      coeffs_in_data_log_force[8018] <= 16'h0000;
      coeffs_in_data_log_force[8019] <= 16'h0000;
      coeffs_in_data_log_force[8020] <= 16'h0000;
      coeffs_in_data_log_force[8021] <= 16'h0000;
      coeffs_in_data_log_force[8022] <= 16'h0000;
      coeffs_in_data_log_force[8023] <= 16'h0000;
      coeffs_in_data_log_force[8024] <= 16'h0000;
      coeffs_in_data_log_force[8025] <= 16'h0000;
      coeffs_in_data_log_force[8026] <= 16'h0000;
      coeffs_in_data_log_force[8027] <= 16'h0000;
      coeffs_in_data_log_force[8028] <= 16'h0000;
      coeffs_in_data_log_force[8029] <= 16'h0000;
      coeffs_in_data_log_force[8030] <= 16'h0000;
      coeffs_in_data_log_force[8031] <= 16'h0000;
      coeffs_in_data_log_force[8032] <= 16'h0000;
      coeffs_in_data_log_force[8033] <= 16'h0000;
      coeffs_in_data_log_force[8034] <= 16'h0000;
      coeffs_in_data_log_force[8035] <= 16'h0000;
      coeffs_in_data_log_force[8036] <= 16'h0000;
      coeffs_in_data_log_force[8037] <= 16'h0000;
      coeffs_in_data_log_force[8038] <= 16'h0000;
      coeffs_in_data_log_force[8039] <= 16'h0000;
      coeffs_in_data_log_force[8040] <= 16'h0000;
      coeffs_in_data_log_force[8041] <= 16'h0000;
      coeffs_in_data_log_force[8042] <= 16'h0000;
      coeffs_in_data_log_force[8043] <= 16'h0000;
      coeffs_in_data_log_force[8044] <= 16'h0000;
      coeffs_in_data_log_force[8045] <= 16'h0000;
      coeffs_in_data_log_force[8046] <= 16'h0000;
      coeffs_in_data_log_force[8047] <= 16'h0000;
      coeffs_in_data_log_force[8048] <= 16'h0000;
      coeffs_in_data_log_force[8049] <= 16'h0000;
      coeffs_in_data_log_force[8050] <= 16'h0000;
      coeffs_in_data_log_force[8051] <= 16'h0000;
      coeffs_in_data_log_force[8052] <= 16'h0000;
      coeffs_in_data_log_force[8053] <= 16'h0000;
      coeffs_in_data_log_force[8054] <= 16'h0000;
      coeffs_in_data_log_force[8055] <= 16'h0000;
      coeffs_in_data_log_force[8056] <= 16'h0000;
      coeffs_in_data_log_force[8057] <= 16'h0000;
      coeffs_in_data_log_force[8058] <= 16'h0000;
      coeffs_in_data_log_force[8059] <= 16'h0000;
      coeffs_in_data_log_force[8060] <= 16'h0000;
      coeffs_in_data_log_force[8061] <= 16'h0000;
      coeffs_in_data_log_force[8062] <= 16'h0000;
      coeffs_in_data_log_force[8063] <= 16'h0000;
      coeffs_in_data_log_force[8064] <= 16'h0000;
      coeffs_in_data_log_force[8065] <= 16'h0000;
      coeffs_in_data_log_force[8066] <= 16'h0000;
      coeffs_in_data_log_force[8067] <= 16'h0000;
      coeffs_in_data_log_force[8068] <= 16'h0000;
      coeffs_in_data_log_force[8069] <= 16'h0000;
      coeffs_in_data_log_force[8070] <= 16'h0000;
      coeffs_in_data_log_force[8071] <= 16'h0000;
      coeffs_in_data_log_force[8072] <= 16'h0000;
      coeffs_in_data_log_force[8073] <= 16'h0000;
      coeffs_in_data_log_force[8074] <= 16'h0000;
      coeffs_in_data_log_force[8075] <= 16'h0000;
      coeffs_in_data_log_force[8076] <= 16'h0000;
      coeffs_in_data_log_force[8077] <= 16'h0000;
      coeffs_in_data_log_force[8078] <= 16'h0000;
      coeffs_in_data_log_force[8079] <= 16'h0000;
      coeffs_in_data_log_force[8080] <= 16'h0000;
      coeffs_in_data_log_force[8081] <= 16'h0000;
      coeffs_in_data_log_force[8082] <= 16'h0000;
      coeffs_in_data_log_force[8083] <= 16'h0000;
      coeffs_in_data_log_force[8084] <= 16'h0000;
      coeffs_in_data_log_force[8085] <= 16'h0000;
      coeffs_in_data_log_force[8086] <= 16'h0000;
      coeffs_in_data_log_force[8087] <= 16'h0000;
      coeffs_in_data_log_force[8088] <= 16'h0000;
      coeffs_in_data_log_force[8089] <= 16'h0000;
      coeffs_in_data_log_force[8090] <= 16'h0000;
      coeffs_in_data_log_force[8091] <= 16'h0000;
      coeffs_in_data_log_force[8092] <= 16'h0000;
      coeffs_in_data_log_force[8093] <= 16'h0000;
      coeffs_in_data_log_force[8094] <= 16'h0000;
      coeffs_in_data_log_force[8095] <= 16'h0000;
      coeffs_in_data_log_force[8096] <= 16'h0000;
      coeffs_in_data_log_force[8097] <= 16'h0000;
      coeffs_in_data_log_force[8098] <= 16'h0000;
      coeffs_in_data_log_force[8099] <= 16'h0000;
      coeffs_in_data_log_force[8100] <= 16'h0000;
      coeffs_in_data_log_force[8101] <= 16'h0000;
      coeffs_in_data_log_force[8102] <= 16'h0000;
      coeffs_in_data_log_force[8103] <= 16'h0000;
      coeffs_in_data_log_force[8104] <= 16'h0000;
      coeffs_in_data_log_force[8105] <= 16'h0000;
      coeffs_in_data_log_force[8106] <= 16'h0000;
      coeffs_in_data_log_force[8107] <= 16'h0000;
      coeffs_in_data_log_force[8108] <= 16'h0000;
      coeffs_in_data_log_force[8109] <= 16'h0000;
      coeffs_in_data_log_force[8110] <= 16'h0000;
      coeffs_in_data_log_force[8111] <= 16'h0000;
      coeffs_in_data_log_force[8112] <= 16'h0000;
      coeffs_in_data_log_force[8113] <= 16'h0000;
      coeffs_in_data_log_force[8114] <= 16'h0000;
      coeffs_in_data_log_force[8115] <= 16'h0000;
      coeffs_in_data_log_force[8116] <= 16'h0000;
      coeffs_in_data_log_force[8117] <= 16'h0000;
      coeffs_in_data_log_force[8118] <= 16'h0000;
      coeffs_in_data_log_force[8119] <= 16'h0000;
      coeffs_in_data_log_force[8120] <= 16'h0000;
      coeffs_in_data_log_force[8121] <= 16'h0000;
      coeffs_in_data_log_force[8122] <= 16'h0000;
      coeffs_in_data_log_force[8123] <= 16'h0000;
      coeffs_in_data_log_force[8124] <= 16'h0000;
      coeffs_in_data_log_force[8125] <= 16'h0000;
      coeffs_in_data_log_force[8126] <= 16'h0000;
      coeffs_in_data_log_force[8127] <= 16'h0000;
      coeffs_in_data_log_force[8128] <= 16'h0000;
      coeffs_in_data_log_force[8129] <= 16'h0000;
      coeffs_in_data_log_force[8130] <= 16'h0000;
      coeffs_in_data_log_force[8131] <= 16'h0000;
      coeffs_in_data_log_force[8132] <= 16'h0000;
      coeffs_in_data_log_force[8133] <= 16'h0000;
      coeffs_in_data_log_force[8134] <= 16'h0000;
      coeffs_in_data_log_force[8135] <= 16'h0000;
      coeffs_in_data_log_force[8136] <= 16'h0000;
      coeffs_in_data_log_force[8137] <= 16'h0000;
      coeffs_in_data_log_force[8138] <= 16'h0000;
      coeffs_in_data_log_force[8139] <= 16'h0000;
      coeffs_in_data_log_force[8140] <= 16'h0000;
      coeffs_in_data_log_force[8141] <= 16'h0000;
      coeffs_in_data_log_force[8142] <= 16'h0000;
      coeffs_in_data_log_force[8143] <= 16'h0000;
      coeffs_in_data_log_force[8144] <= 16'h0000;
      coeffs_in_data_log_force[8145] <= 16'h0000;
      coeffs_in_data_log_force[8146] <= 16'h0000;
      coeffs_in_data_log_force[8147] <= 16'h0000;
      coeffs_in_data_log_force[8148] <= 16'h0000;
      coeffs_in_data_log_force[8149] <= 16'h0000;
      coeffs_in_data_log_force[8150] <= 16'h0000;
      coeffs_in_data_log_force[8151] <= 16'h0000;
      coeffs_in_data_log_force[8152] <= 16'h0000;
      coeffs_in_data_log_force[8153] <= 16'h0000;
      coeffs_in_data_log_force[8154] <= 16'h0000;
      coeffs_in_data_log_force[8155] <= 16'h0000;
      coeffs_in_data_log_force[8156] <= 16'h0000;
      coeffs_in_data_log_force[8157] <= 16'h0000;
      coeffs_in_data_log_force[8158] <= 16'h0000;
      coeffs_in_data_log_force[8159] <= 16'h0000;
      coeffs_in_data_log_force[8160] <= 16'h0000;
      coeffs_in_data_log_force[8161] <= 16'h0000;
      coeffs_in_data_log_force[8162] <= 16'h0000;
      coeffs_in_data_log_force[8163] <= 16'h0000;
      coeffs_in_data_log_force[8164] <= 16'h0000;
      coeffs_in_data_log_force[8165] <= 16'h0000;
      coeffs_in_data_log_force[8166] <= 16'h0000;
      coeffs_in_data_log_force[8167] <= 16'h0000;
      coeffs_in_data_log_force[8168] <= 16'h0000;
      coeffs_in_data_log_force[8169] <= 16'h0000;
      coeffs_in_data_log_force[8170] <= 16'h0000;
      coeffs_in_data_log_force[8171] <= 16'h0000;
      coeffs_in_data_log_force[8172] <= 16'h0000;
      coeffs_in_data_log_force[8173] <= 16'h0000;
      coeffs_in_data_log_force[8174] <= 16'h0000;
      coeffs_in_data_log_force[8175] <= 16'h0000;
      coeffs_in_data_log_force[8176] <= 16'h0000;
      coeffs_in_data_log_force[8177] <= 16'h0000;
      coeffs_in_data_log_force[8178] <= 16'h0000;
      coeffs_in_data_log_force[8179] <= 16'h0000;
      coeffs_in_data_log_force[8180] <= 16'h0000;
      coeffs_in_data_log_force[8181] <= 16'h0000;
      coeffs_in_data_log_force[8182] <= 16'h0000;
      coeffs_in_data_log_force[8183] <= 16'h0000;
      coeffs_in_data_log_force[8184] <= 16'h0000;
      coeffs_in_data_log_force[8185] <= 16'h0000;
      coeffs_in_data_log_force[8186] <= 16'h0000;
      coeffs_in_data_log_force[8187] <= 16'h0000;
      coeffs_in_data_log_force[8188] <= 16'h0000;
      coeffs_in_data_log_force[8189] <= 16'h0000;
      coeffs_in_data_log_force[8190] <= 16'h0000;
      coeffs_in_data_log_force[8191] <= 16'h0000;
      coeffs_in_data_log_force[8192] <= 16'h0000;
      coeffs_in_data_log_force[8193] <= 16'h0000;
      coeffs_in_data_log_force[8194] <= 16'h0000;
      coeffs_in_data_log_force[8195] <= 16'h0000;
      coeffs_in_data_log_force[8196] <= 16'h0000;
      coeffs_in_data_log_force[8197] <= 16'h0000;
      coeffs_in_data_log_force[8198] <= 16'h0000;
      coeffs_in_data_log_force[8199] <= 16'h0000;
      coeffs_in_data_log_force[8200] <= 16'h0000;
      coeffs_in_data_log_force[8201] <= 16'h0000;
      coeffs_in_data_log_force[8202] <= 16'h0000;
      coeffs_in_data_log_force[8203] <= 16'h0000;
      coeffs_in_data_log_force[8204] <= 16'h0000;
      coeffs_in_data_log_force[8205] <= 16'h0000;
      coeffs_in_data_log_force[8206] <= 16'h0000;
      coeffs_in_data_log_force[8207] <= 16'h0000;
      coeffs_in_data_log_force[8208] <= 16'h0000;
      coeffs_in_data_log_force[8209] <= 16'h0000;
      coeffs_in_data_log_force[8210] <= 16'h0000;
      coeffs_in_data_log_force[8211] <= 16'h0000;
      coeffs_in_data_log_force[8212] <= 16'h0000;
      coeffs_in_data_log_force[8213] <= 16'h0000;
      coeffs_in_data_log_force[8214] <= 16'h0000;
      coeffs_in_data_log_force[8215] <= 16'h0000;
      coeffs_in_data_log_force[8216] <= 16'h0000;
      coeffs_in_data_log_force[8217] <= 16'h0000;
      coeffs_in_data_log_force[8218] <= 16'h0000;
      coeffs_in_data_log_force[8219] <= 16'h0000;
      coeffs_in_data_log_force[8220] <= 16'h0000;
      coeffs_in_data_log_force[8221] <= 16'h0000;
      coeffs_in_data_log_force[8222] <= 16'h0000;
      coeffs_in_data_log_force[8223] <= 16'h0000;
      coeffs_in_data_log_force[8224] <= 16'h0000;
      coeffs_in_data_log_force[8225] <= 16'h0000;
      coeffs_in_data_log_force[8226] <= 16'h0000;
      coeffs_in_data_log_force[8227] <= 16'h0000;
      coeffs_in_data_log_force[8228] <= 16'h0000;
      coeffs_in_data_log_force[8229] <= 16'h0000;
      coeffs_in_data_log_force[8230] <= 16'h0000;
      coeffs_in_data_log_force[8231] <= 16'h0000;
      coeffs_in_data_log_force[8232] <= 16'h0000;
      coeffs_in_data_log_force[8233] <= 16'h0000;
      coeffs_in_data_log_force[8234] <= 16'h0000;
      coeffs_in_data_log_force[8235] <= 16'h0000;
      coeffs_in_data_log_force[8236] <= 16'h0000;
      coeffs_in_data_log_force[8237] <= 16'h0000;
      coeffs_in_data_log_force[8238] <= 16'h0000;
      coeffs_in_data_log_force[8239] <= 16'h0000;
      coeffs_in_data_log_force[8240] <= 16'h0000;
      coeffs_in_data_log_force[8241] <= 16'h0000;
      coeffs_in_data_log_force[8242] <= 16'h0000;
      coeffs_in_data_log_force[8243] <= 16'h0000;
      coeffs_in_data_log_force[8244] <= 16'h0000;
      coeffs_in_data_log_force[8245] <= 16'h0000;
      coeffs_in_data_log_force[8246] <= 16'h0000;
      coeffs_in_data_log_force[8247] <= 16'h0000;
      coeffs_in_data_log_force[8248] <= 16'h0000;
      coeffs_in_data_log_force[8249] <= 16'h0000;
      coeffs_in_data_log_force[8250] <= 16'h0000;
      coeffs_in_data_log_force[8251] <= 16'h0000;
      coeffs_in_data_log_force[8252] <= 16'h0000;
      coeffs_in_data_log_force[8253] <= 16'h0000;
      coeffs_in_data_log_force[8254] <= 16'h0000;
      coeffs_in_data_log_force[8255] <= 16'h0000;
      coeffs_in_data_log_force[8256] <= 16'h0000;
      coeffs_in_data_log_force[8257] <= 16'h0000;
      coeffs_in_data_log_force[8258] <= 16'h0000;
      coeffs_in_data_log_force[8259] <= 16'h0000;
      coeffs_in_data_log_force[8260] <= 16'h0000;
      coeffs_in_data_log_force[8261] <= 16'h0000;
      coeffs_in_data_log_force[8262] <= 16'h0000;
      coeffs_in_data_log_force[8263] <= 16'h0000;
      coeffs_in_data_log_force[8264] <= 16'h0000;
      coeffs_in_data_log_force[8265] <= 16'h0000;
      coeffs_in_data_log_force[8266] <= 16'h0000;
      coeffs_in_data_log_force[8267] <= 16'h0000;
      coeffs_in_data_log_force[8268] <= 16'h0000;
      coeffs_in_data_log_force[8269] <= 16'h0000;
      coeffs_in_data_log_force[8270] <= 16'h0000;
      coeffs_in_data_log_force[8271] <= 16'h0000;
      coeffs_in_data_log_force[8272] <= 16'h0000;
      coeffs_in_data_log_force[8273] <= 16'h0000;
      coeffs_in_data_log_force[8274] <= 16'h0000;
      coeffs_in_data_log_force[8275] <= 16'h0000;
      coeffs_in_data_log_force[8276] <= 16'h0000;
      coeffs_in_data_log_force[8277] <= 16'h0000;
      coeffs_in_data_log_force[8278] <= 16'h0000;
      coeffs_in_data_log_force[8279] <= 16'h0000;
      coeffs_in_data_log_force[8280] <= 16'h0000;
      coeffs_in_data_log_force[8281] <= 16'h0000;
      coeffs_in_data_log_force[8282] <= 16'h0000;
      coeffs_in_data_log_force[8283] <= 16'h0000;
      coeffs_in_data_log_force[8284] <= 16'h0000;
      coeffs_in_data_log_force[8285] <= 16'h0000;
      coeffs_in_data_log_force[8286] <= 16'h0000;
      coeffs_in_data_log_force[8287] <= 16'h0000;
      coeffs_in_data_log_force[8288] <= 16'h0000;
      coeffs_in_data_log_force[8289] <= 16'h0000;
      coeffs_in_data_log_force[8290] <= 16'h0000;
      coeffs_in_data_log_force[8291] <= 16'h0000;
      coeffs_in_data_log_force[8292] <= 16'h0000;
      coeffs_in_data_log_force[8293] <= 16'h0000;
      coeffs_in_data_log_force[8294] <= 16'h0000;
      coeffs_in_data_log_force[8295] <= 16'h0000;
      coeffs_in_data_log_force[8296] <= 16'h0000;
      coeffs_in_data_log_force[8297] <= 16'h0000;
      coeffs_in_data_log_force[8298] <= 16'h0000;
      coeffs_in_data_log_force[8299] <= 16'h0000;
      coeffs_in_data_log_force[8300] <= 16'h0000;
      coeffs_in_data_log_force[8301] <= 16'h0000;
      coeffs_in_data_log_force[8302] <= 16'h0000;
      coeffs_in_data_log_force[8303] <= 16'h0000;
      coeffs_in_data_log_force[8304] <= 16'h0000;
      coeffs_in_data_log_force[8305] <= 16'h0000;
      coeffs_in_data_log_force[8306] <= 16'h0000;
      coeffs_in_data_log_force[8307] <= 16'h0000;
      coeffs_in_data_log_force[8308] <= 16'h0000;
      coeffs_in_data_log_force[8309] <= 16'h0000;
      coeffs_in_data_log_force[8310] <= 16'h0000;
      coeffs_in_data_log_force[8311] <= 16'h0000;
      coeffs_in_data_log_force[8312] <= 16'h0000;
      coeffs_in_data_log_force[8313] <= 16'h0000;
      coeffs_in_data_log_force[8314] <= 16'h0000;
      coeffs_in_data_log_force[8315] <= 16'h0000;
      coeffs_in_data_log_force[8316] <= 16'h0000;
      coeffs_in_data_log_force[8317] <= 16'h0000;
      coeffs_in_data_log_force[8318] <= 16'h0000;
      coeffs_in_data_log_force[8319] <= 16'h0000;

      // Output data for filter_out
      filter_out_expected[  0] <= 16'h0000;
      filter_out_expected[  1] <= 16'h0000;
      filter_out_expected[  2] <= 16'hffff;
      filter_out_expected[  3] <= 16'hffff;
      filter_out_expected[  4] <= 16'hffff;
      filter_out_expected[  5] <= 16'hffff;
      filter_out_expected[  6] <= 16'hffff;
      filter_out_expected[  7] <= 16'hffff;
      filter_out_expected[  8] <= 16'hffff;
      filter_out_expected[  9] <= 16'hffff;
      filter_out_expected[ 10] <= 16'h0000;
      filter_out_expected[ 11] <= 16'h0000;
      filter_out_expected[ 12] <= 16'h0000;
      filter_out_expected[ 13] <= 16'h0000;
      filter_out_expected[ 14] <= 16'h0000;
      filter_out_expected[ 15] <= 16'h0000;
      filter_out_expected[ 16] <= 16'h0000;
      filter_out_expected[ 17] <= 16'h0000;
      filter_out_expected[ 18] <= 16'hffff;
      filter_out_expected[ 19] <= 16'hffff;
      filter_out_expected[ 20] <= 16'hffff;
      filter_out_expected[ 21] <= 16'hffff;
      filter_out_expected[ 22] <= 16'hffff;
      filter_out_expected[ 23] <= 16'hffff;
      filter_out_expected[ 24] <= 16'hffff;
      filter_out_expected[ 25] <= 16'hffff;
      filter_out_expected[ 26] <= 16'h0000;
      filter_out_expected[ 27] <= 16'h0000;
      filter_out_expected[ 28] <= 16'h0000;
      filter_out_expected[ 29] <= 16'h0000;
      filter_out_expected[ 30] <= 16'h0000;
      filter_out_expected[ 31] <= 16'h0000;
      filter_out_expected[ 32] <= 16'h0000;
      filter_out_expected[ 33] <= 16'h0000;
      filter_out_expected[ 34] <= 16'h0000;
      filter_out_expected[ 35] <= 16'h0000;
      filter_out_expected[ 36] <= 16'h0000;
      filter_out_expected[ 37] <= 16'h0000;
      filter_out_expected[ 38] <= 16'h0000;
      filter_out_expected[ 39] <= 16'h0000;
      filter_out_expected[ 40] <= 16'h0000;
      filter_out_expected[ 41] <= 16'h0000;
      filter_out_expected[ 42] <= 16'hffff;
      filter_out_expected[ 43] <= 16'hffff;
      filter_out_expected[ 44] <= 16'hffff;
      filter_out_expected[ 45] <= 16'hffff;
      filter_out_expected[ 46] <= 16'hffff;
      filter_out_expected[ 47] <= 16'hffff;
      filter_out_expected[ 48] <= 16'hffff;
      filter_out_expected[ 49] <= 16'hffff;
      filter_out_expected[ 50] <= 16'h0000;
      filter_out_expected[ 51] <= 16'h0000;
      filter_out_expected[ 52] <= 16'h0000;
      filter_out_expected[ 53] <= 16'h0000;
      filter_out_expected[ 54] <= 16'h0000;
      filter_out_expected[ 55] <= 16'h0000;
      filter_out_expected[ 56] <= 16'h0000;
      filter_out_expected[ 57] <= 16'h0000;
      filter_out_expected[ 58] <= 16'hffff;
      filter_out_expected[ 59] <= 16'hffff;
      filter_out_expected[ 60] <= 16'hffff;
      filter_out_expected[ 61] <= 16'hffff;
      filter_out_expected[ 62] <= 16'hffff;
      filter_out_expected[ 63] <= 16'hffff;
      filter_out_expected[ 64] <= 16'hffff;
      filter_out_expected[ 65] <= 16'hffff;
      filter_out_expected[ 66] <= 16'h0000;
      filter_out_expected[ 67] <= 16'h0000;
      filter_out_expected[ 68] <= 16'h0000;
      filter_out_expected[ 69] <= 16'h0000;
      filter_out_expected[ 70] <= 16'h0000;
      filter_out_expected[ 71] <= 16'h0000;
      filter_out_expected[ 72] <= 16'h0000;
      filter_out_expected[ 73] <= 16'h0000;
      filter_out_expected[ 74] <= 16'h0000;
      filter_out_expected[ 75] <= 16'h0000;
      filter_out_expected[ 76] <= 16'h0000;
      filter_out_expected[ 77] <= 16'h0000;
      filter_out_expected[ 78] <= 16'h0000;
      filter_out_expected[ 79] <= 16'h0000;
      filter_out_expected[ 80] <= 16'h0000;
      filter_out_expected[ 81] <= 16'h0000;
      filter_out_expected[ 82] <= 16'h0000;
      filter_out_expected[ 83] <= 16'h0000;
      filter_out_expected[ 84] <= 16'h0000;
      filter_out_expected[ 85] <= 16'h0000;
      filter_out_expected[ 86] <= 16'h0000;
      filter_out_expected[ 87] <= 16'h0000;
      filter_out_expected[ 88] <= 16'h0000;
      filter_out_expected[ 89] <= 16'h0000;
      filter_out_expected[ 90] <= 16'h0000;
      filter_out_expected[ 91] <= 16'h0000;
      filter_out_expected[ 92] <= 16'h0000;
      filter_out_expected[ 93] <= 16'h0000;
      filter_out_expected[ 94] <= 16'h0000;
      filter_out_expected[ 95] <= 16'h0000;
      filter_out_expected[ 96] <= 16'h0000;
      filter_out_expected[ 97] <= 16'h0000;
      filter_out_expected[ 98] <= 16'h0000;
      filter_out_expected[ 99] <= 16'h0000;
      filter_out_expected[100] <= 16'h0000;
      filter_out_expected[101] <= 16'h0000;
      filter_out_expected[102] <= 16'h0000;
      filter_out_expected[103] <= 16'h0000;
      filter_out_expected[104] <= 16'h0000;
      filter_out_expected[105] <= 16'h0000;
      filter_out_expected[106] <= 16'h0000;
      filter_out_expected[107] <= 16'h0000;
      filter_out_expected[108] <= 16'h0000;
      filter_out_expected[109] <= 16'h0000;
      filter_out_expected[110] <= 16'h0000;
      filter_out_expected[111] <= 16'h0000;
      filter_out_expected[112] <= 16'h0000;
      filter_out_expected[113] <= 16'h0000;
      filter_out_expected[114] <= 16'h0000;
      filter_out_expected[115] <= 16'h0000;
      filter_out_expected[116] <= 16'h0000;
      filter_out_expected[117] <= 16'h0000;
      filter_out_expected[118] <= 16'h0000;
      filter_out_expected[119] <= 16'h0000;
      filter_out_expected[120] <= 16'h0000;
      filter_out_expected[121] <= 16'h0000;
      filter_out_expected[122] <= 16'h0000;
      filter_out_expected[123] <= 16'h0000;
      filter_out_expected[124] <= 16'h0000;
      filter_out_expected[125] <= 16'h0000;
      filter_out_expected[126] <= 16'h0000;
      filter_out_expected[127] <= 16'h0000;
      filter_out_expected[128] <= 16'h0000;
      filter_out_expected[129] <= 16'h0000;

    end  // Input & Output data
  //************************************


  parameter MAX_ERROR_COUNT = 130;  //uint32


  // Signals
  reg clk;  // boolean
  reg clk_enable;  // boolean
  reg rst;  // boolean
  reg signed [15:0] filter_in;  // sfix16
  reg write_enable;  // boolean
  reg write_done;  // boolean
  reg [5:0] write_address;  // ufix6
  reg signed [15:0] coeffs_in;  // sfix16_En18
  wire signed [15:0] filter_out;  // sfix16

  reg tb_enb;  // boolean
  wire srcDone;  // boolean
  wire snkDone;  // boolean
  wire testFailure;  // boolean
  reg tbenb_dly;  // boolean
  reg [5:0] counter;  // ufix6
  wire phase_1;  // boolean
  wire phase_all;  // boolean
  wire phase_all_1;  // boolean
  wire phase_all_2;  // boolean
  wire phase_all_3;  // boolean
  wire rdEnb_phase_1;  // boolean
  wire rdEnb_phase_all;  // boolean
  wire filter_in_data_log_rdenb;  // boolean
  reg [7:0] filter_in_data_log_addr;  // ufix8
  reg filter_in_data_log_done;  // boolean
  wire signed [15:0] rawData_filter_in;  // sfix16
  reg signed [15:0] holdData_filter_in;  // sfix16
  wire write_enable_data_log_rdenb;  // boolean
  reg [13:0] write_enable_data_log_addr;  // ufix14
  reg write_enable_data_log_done;  // boolean
  wire rawData_write_enable;  // boolean
  reg holdData_write_enable;  // boolean
  wire write_done_data_log_rdenb;  // boolean
  reg [13:0] write_done_data_log_addr;  // ufix14
  reg write_done_data_log_done;  // boolean
  wire rawData_write_done;  // boolean
  reg holdData_write_done;  // boolean
  wire write_address_data_log_rdenb;  // boolean
  reg [13:0] write_address_data_log_addr;  // ufix14
  reg write_address_data_log_done;  // boolean
  wire [5:0] rawData_write_address;  // ufix6
  reg [5:0] holdData_write_address;  // ufix6
  wire coeffs_in_data_log_rdenb;  // boolean
  reg [13:0] coeffs_in_data_log_addr;  // ufix14
  reg coeffs_in_data_log_done;  // boolean
  wire signed [15:0] rawData_coeffs_in;  // sfix16_En18
  reg signed [15:0] holdData_coeffs_in;  // sfix16_En18
  reg filter_out_testFailure;  // boolean
  integer filter_out_errCnt;  // uint32
  wire delayLine_out;  // boolean
  wire expected_ce_out;  // boolean
  reg int_delay_pipe[0:128];  // boolean
  wire filter_out_rdenb;  // boolean
  reg [7:0] filter_out_addr;  // ufix8
  reg filter_out_done;  // boolean
  wire signed [15:0] filter_out_ref;  // sfix16
  wire signed [15:0] filter_out_dataTable;  // sfix16
  wire signed [15:0] filter_out_refTmp;  // sfix16
  reg signed [15:0] regout;  // sfix16
  reg check1_Done;  // boolean

  // Module Instances
  filter u_filter (
      .clk(clk),
      .clk_enable(clk_enable),
      .rst(rst),
      .filter_in(filter_in),
      .write_enable(write_enable),
      .write_done(write_done),
      .write_address(write_address),
      .coeffs_in(coeffs_in),
      .filter_out(filter_out)
  );


  // Block Statements
  // -------------------------------------------------------------
  // Driving the test bench enable
  // -------------------------------------------------------------

  always @(rst, snkDone) begin
    if (rst == 1'b1) tb_enb <= 1'b0;
    else if (snkDone == 1'b0) tb_enb <= 1'b1;
    else begin
      #(clk_period * 2);
      tb_enb <= 1'b0;
    end
  end

  always @(posedge clk or posedge rst) // completed_msg
  begin
    if (rst) begin
      // Nothing to reset.
    end else begin
      if (snkDone == 1) begin
        if (testFailure == 0) $display("**************TEST COMPLETED (PASSED)**************");
        else $display("**************TEST COMPLETED (FAILED)**************");
      end
    end
  end  // completed_msg;

  // -------------------------------------------------------------
  // System Clock (fast clock) and reset
  // -------------------------------------------------------------

  always  // clock generation
  begin // clk_gen
    clk <= 1'b1;
    #clk_high;
    clk <= 1'b0;
    #clk_low;
    if (snkDone == 1) begin
      clk <= 1'b1;
      #clk_high;
      clk <= 1'b0;
      #clk_low;
      $stop;
    end
  end  // clk_gen

  initial  // reset block
    begin  // rst_gen
      rst <= 1'b1;
      #(clk_period * 2);
      @(posedge clk);
      #(clk_hold);
      rst <= 1'b0;
    end  // rst_gen

  // -------------------------------------------------------------
  // Testbench clock enable
  // -------------------------------------------------------------

  always @(posedge clk or posedge rst) begin : tb_enb_delay
    if (rst == 1'b1) begin
      tbenb_dly <= 1'b0;
    end else begin
      if (tb_enb == 1'b1) begin
        tbenb_dly <= tb_enb;
      end
    end
  end  // tb_enb_delay

  // -------------------------------------------------------------
  // Slow Clock (clkenb)
  // -------------------------------------------------------------

  always @(posedge clk or posedge rst) begin : slow_clock_enable
    if (rst == 1'b1) begin
      counter <= 6'b000001;
    end else begin
      if (tbenb_dly == 1'b1) begin
        if (counter >= 6'b111111) begin
          counter <= 6'b000000;
        end else begin
          counter <= counter + 6'b000001;
        end
      end
    end
  end  // slow_clock_enable

  assign phase_1 = (counter == 6'b000001 && tbenb_dly == 1'b1) ? 1'b1 : 1'b0;

  assign phase_all = tbenb_dly ? 1'b1 : 1'b0;

  assign phase_all_1 = tbenb_dly ? 1'b1 : 1'b0;

  assign phase_all_2 = tbenb_dly ? 1'b1 : 1'b0;

  assign phase_all_3 = tbenb_dly ? 1'b1 : 1'b0;

  assign rdEnb_phase_1 = phase_1;

  assign rdEnb_phase_all = phase_all;

  // -------------------------------------------------------------
  // Read the data and transmit it to the DUT
  // -------------------------------------------------------------

  always @(posedge clk or posedge rst) begin
    filter_in_data_log_task(clk, rst, filter_in_data_log_rdenb, filter_in_data_log_addr,
                            filter_in_data_log_done);
  end

  assign filter_in_data_log_rdenb = rdEnb_phase_1;

  assign rawData_filter_in = filter_in_data_log_force[filter_in_data_log_addr];

  always @(posedge clk or posedge rst) begin  // stimuli_filter_in_data_log_filter_in_reg
    if (rst) begin
      holdData_filter_in <= 16'b0;
    end else begin
      holdData_filter_in <= rawData_filter_in;
    end
  end

  always @ (filter_in_data_log_rdenb, filter_in_data_log_addr, tbenb_dly)
  begin // stimuli_filter_in_data_log_filter_in
    if (tbenb_dly == 0) begin
      filter_in <= #clk_hold 16'b0;
    end else if (filter_in_data_log_rdenb == 1) begin
      filter_in <= #clk_hold rawData_filter_in;
    end else begin
      filter_in <= #clk_hold holdData_filter_in;
    end
  end  // stimuli_filter_in_data_log_filter_in

  // -------------------------------------------------------------
  // Read the data and transmit it to the DUT
  // -------------------------------------------------------------

  always @(posedge clk or posedge rst) begin
    write_enable_data_log_task(clk, rst, write_enable_data_log_rdenb, write_enable_data_log_addr,
                               write_enable_data_log_done);
  end

  assign write_enable_data_log_rdenb = rdEnb_phase_all;

  assign rawData_write_enable = write_enable_data_log_force[write_enable_data_log_addr];

  always @(posedge clk or posedge rst) begin  // stimuli_write_enable_data_log_write_enable_reg
    if (rst) begin
      holdData_write_enable <= 1'b0;
    end else begin
      holdData_write_enable <= rawData_write_enable;
    end
  end

  always @ (write_enable_data_log_rdenb, write_enable_data_log_addr, tbenb_dly)
  begin // stimuli_write_enable_data_log_write_enable
    if (tbenb_dly == 0) begin
      write_enable <= #clk_hold 1'b0;
    end else if (write_enable_data_log_rdenb == 1) begin
      write_enable <= #clk_hold rawData_write_enable;
    end else begin
      write_enable <= #clk_hold holdData_write_enable;
    end
  end  // stimuli_write_enable_data_log_write_enable

  // -------------------------------------------------------------
  // Read the data and transmit it to the DUT
  // -------------------------------------------------------------

  always @(posedge clk or posedge rst) begin
    write_done_data_log_task(clk, rst, write_done_data_log_rdenb, write_done_data_log_addr,
                             write_done_data_log_done);
  end

  assign write_done_data_log_rdenb = rdEnb_phase_all;

  assign rawData_write_done = write_done_data_log_force[write_done_data_log_addr];

  always @(posedge clk or posedge rst) begin  // stimuli_write_done_data_log_write_done_reg
    if (rst) begin
      holdData_write_done <= 1'b0;
    end else begin
      holdData_write_done <= rawData_write_done;
    end
  end

  always @ (write_done_data_log_rdenb, write_done_data_log_addr, tbenb_dly)
  begin // stimuli_write_done_data_log_write_done
    if (tbenb_dly == 0) begin
      write_done <= #clk_hold 1'b0;
    end else if (write_done_data_log_rdenb == 1) begin
      write_done <= #clk_hold rawData_write_done;
    end else begin
      write_done <= #clk_hold holdData_write_done;
    end
  end  // stimuli_write_done_data_log_write_done

  // -------------------------------------------------------------
  // Read the data and transmit it to the DUT
  // -------------------------------------------------------------

  always @(posedge clk or posedge rst) begin
    write_address_data_log_task(clk, rst, write_address_data_log_rdenb, write_address_data_log_addr,
                                write_address_data_log_done);
  end

  assign write_address_data_log_rdenb = rdEnb_phase_all;

  assign rawData_write_address = write_address_data_log_force[write_address_data_log_addr];

  always @(posedge clk or posedge rst) begin  // stimuli_write_address_data_log_write_address_reg
    if (rst) begin
      holdData_write_address <= 6'b0;
    end else begin
      holdData_write_address <= rawData_write_address;
    end
  end

  always @ (write_address_data_log_rdenb, write_address_data_log_addr, tbenb_dly)
  begin // stimuli_write_address_data_log_write_address
    if (tbenb_dly == 0) begin
      write_address <= #clk_hold 6'b0;
    end else if (write_address_data_log_rdenb == 1) begin
      write_address <= #clk_hold rawData_write_address;
    end else begin
      write_address <= #clk_hold holdData_write_address;
    end
  end  // stimuli_write_address_data_log_write_address

  // -------------------------------------------------------------
  // Read the data and transmit it to the DUT
  // -------------------------------------------------------------

  always @(posedge clk or posedge rst) begin
    coeffs_in_data_log_task(clk, rst, coeffs_in_data_log_rdenb, coeffs_in_data_log_addr,
                            coeffs_in_data_log_done);
  end

  assign coeffs_in_data_log_rdenb = rdEnb_phase_all;

  assign rawData_coeffs_in = coeffs_in_data_log_force[coeffs_in_data_log_addr];

  always @(posedge clk or posedge rst) begin  // stimuli_coeffs_in_data_log_coeffs_in_reg
    if (rst) begin
      holdData_coeffs_in <= 18'b0;
    end else begin
      holdData_coeffs_in <= rawData_coeffs_in;
    end
  end

  always @ (coeffs_in_data_log_rdenb, coeffs_in_data_log_addr, tbenb_dly)
  begin // stimuli_coeffs_in_data_log_coeffs_in
    if (tbenb_dly == 0) begin
      coeffs_in <= #clk_hold 18'b0;
    end else if (coeffs_in_data_log_rdenb == 1) begin
      coeffs_in <= #clk_hold rawData_coeffs_in;
    end else begin
      coeffs_in <= #clk_hold holdData_coeffs_in;
    end
  end  // stimuli_coeffs_in_data_log_coeffs_in

  // -------------------------------------------------------------
  // Create done signal for Input data
  // -------------------------------------------------------------

  assign srcDone = filter_in_data_log_done && write_enable_data_log_done && write_done_data_log_done && write_address_data_log_done && coeffs_in_data_log_done;


  always @(posedge clk or posedge rst) begin : ceout_delayLine
    if (rst == 1'b1) begin
      int_delay_pipe[0]   <= 1'b0;
      int_delay_pipe[1]   <= 1'b0;
      int_delay_pipe[2]   <= 1'b0;
      int_delay_pipe[3]   <= 1'b0;
      int_delay_pipe[4]   <= 1'b0;
      int_delay_pipe[5]   <= 1'b0;
      int_delay_pipe[6]   <= 1'b0;
      int_delay_pipe[7]   <= 1'b0;
      int_delay_pipe[8]   <= 1'b0;
      int_delay_pipe[9]   <= 1'b0;
      int_delay_pipe[10]  <= 1'b0;
      int_delay_pipe[11]  <= 1'b0;
      int_delay_pipe[12]  <= 1'b0;
      int_delay_pipe[13]  <= 1'b0;
      int_delay_pipe[14]  <= 1'b0;
      int_delay_pipe[15]  <= 1'b0;
      int_delay_pipe[16]  <= 1'b0;
      int_delay_pipe[17]  <= 1'b0;
      int_delay_pipe[18]  <= 1'b0;
      int_delay_pipe[19]  <= 1'b0;
      int_delay_pipe[20]  <= 1'b0;
      int_delay_pipe[21]  <= 1'b0;
      int_delay_pipe[22]  <= 1'b0;
      int_delay_pipe[23]  <= 1'b0;
      int_delay_pipe[24]  <= 1'b0;
      int_delay_pipe[25]  <= 1'b0;
      int_delay_pipe[26]  <= 1'b0;
      int_delay_pipe[27]  <= 1'b0;
      int_delay_pipe[28]  <= 1'b0;
      int_delay_pipe[29]  <= 1'b0;
      int_delay_pipe[30]  <= 1'b0;
      int_delay_pipe[31]  <= 1'b0;
      int_delay_pipe[32]  <= 1'b0;
      int_delay_pipe[33]  <= 1'b0;
      int_delay_pipe[34]  <= 1'b0;
      int_delay_pipe[35]  <= 1'b0;
      int_delay_pipe[36]  <= 1'b0;
      int_delay_pipe[37]  <= 1'b0;
      int_delay_pipe[38]  <= 1'b0;
      int_delay_pipe[39]  <= 1'b0;
      int_delay_pipe[40]  <= 1'b0;
      int_delay_pipe[41]  <= 1'b0;
      int_delay_pipe[42]  <= 1'b0;
      int_delay_pipe[43]  <= 1'b0;
      int_delay_pipe[44]  <= 1'b0;
      int_delay_pipe[45]  <= 1'b0;
      int_delay_pipe[46]  <= 1'b0;
      int_delay_pipe[47]  <= 1'b0;
      int_delay_pipe[48]  <= 1'b0;
      int_delay_pipe[49]  <= 1'b0;
      int_delay_pipe[50]  <= 1'b0;
      int_delay_pipe[51]  <= 1'b0;
      int_delay_pipe[52]  <= 1'b0;
      int_delay_pipe[53]  <= 1'b0;
      int_delay_pipe[54]  <= 1'b0;
      int_delay_pipe[55]  <= 1'b0;
      int_delay_pipe[56]  <= 1'b0;
      int_delay_pipe[57]  <= 1'b0;
      int_delay_pipe[58]  <= 1'b0;
      int_delay_pipe[59]  <= 1'b0;
      int_delay_pipe[60]  <= 1'b0;
      int_delay_pipe[61]  <= 1'b0;
      int_delay_pipe[62]  <= 1'b0;
      int_delay_pipe[63]  <= 1'b0;
      int_delay_pipe[64]  <= 1'b0;
      int_delay_pipe[65]  <= 1'b0;
      int_delay_pipe[66]  <= 1'b0;
      int_delay_pipe[67]  <= 1'b0;
      int_delay_pipe[68]  <= 1'b0;
      int_delay_pipe[69]  <= 1'b0;
      int_delay_pipe[70]  <= 1'b0;
      int_delay_pipe[71]  <= 1'b0;
      int_delay_pipe[72]  <= 1'b0;
      int_delay_pipe[73]  <= 1'b0;
      int_delay_pipe[74]  <= 1'b0;
      int_delay_pipe[75]  <= 1'b0;
      int_delay_pipe[76]  <= 1'b0;
      int_delay_pipe[77]  <= 1'b0;
      int_delay_pipe[78]  <= 1'b0;
      int_delay_pipe[79]  <= 1'b0;
      int_delay_pipe[80]  <= 1'b0;
      int_delay_pipe[81]  <= 1'b0;
      int_delay_pipe[82]  <= 1'b0;
      int_delay_pipe[83]  <= 1'b0;
      int_delay_pipe[84]  <= 1'b0;
      int_delay_pipe[85]  <= 1'b0;
      int_delay_pipe[86]  <= 1'b0;
      int_delay_pipe[87]  <= 1'b0;
      int_delay_pipe[88]  <= 1'b0;
      int_delay_pipe[89]  <= 1'b0;
      int_delay_pipe[90]  <= 1'b0;
      int_delay_pipe[91]  <= 1'b0;
      int_delay_pipe[92]  <= 1'b0;
      int_delay_pipe[93]  <= 1'b0;
      int_delay_pipe[94]  <= 1'b0;
      int_delay_pipe[95]  <= 1'b0;
      int_delay_pipe[96]  <= 1'b0;
      int_delay_pipe[97]  <= 1'b0;
      int_delay_pipe[98]  <= 1'b0;
      int_delay_pipe[99]  <= 1'b0;
      int_delay_pipe[100] <= 1'b0;
      int_delay_pipe[101] <= 1'b0;
      int_delay_pipe[102] <= 1'b0;
      int_delay_pipe[103] <= 1'b0;
      int_delay_pipe[104] <= 1'b0;
      int_delay_pipe[105] <= 1'b0;
      int_delay_pipe[106] <= 1'b0;
      int_delay_pipe[107] <= 1'b0;
      int_delay_pipe[108] <= 1'b0;
      int_delay_pipe[109] <= 1'b0;
      int_delay_pipe[110] <= 1'b0;
      int_delay_pipe[111] <= 1'b0;
      int_delay_pipe[112] <= 1'b0;
      int_delay_pipe[113] <= 1'b0;
      int_delay_pipe[114] <= 1'b0;
      int_delay_pipe[115] <= 1'b0;
      int_delay_pipe[116] <= 1'b0;
      int_delay_pipe[117] <= 1'b0;
      int_delay_pipe[118] <= 1'b0;
      int_delay_pipe[119] <= 1'b0;
      int_delay_pipe[120] <= 1'b0;
      int_delay_pipe[121] <= 1'b0;
      int_delay_pipe[122] <= 1'b0;
      int_delay_pipe[123] <= 1'b0;
      int_delay_pipe[124] <= 1'b0;
      int_delay_pipe[125] <= 1'b0;
      int_delay_pipe[126] <= 1'b0;
      int_delay_pipe[127] <= 1'b0;
      int_delay_pipe[128] <= 1'b0;
    end else begin
      if (clk_enable == 1'b1) begin
        int_delay_pipe[0]   <= rdEnb_phase_1;
        int_delay_pipe[1]   <= int_delay_pipe[0];
        int_delay_pipe[2]   <= int_delay_pipe[1];
        int_delay_pipe[3]   <= int_delay_pipe[2];
        int_delay_pipe[4]   <= int_delay_pipe[3];
        int_delay_pipe[5]   <= int_delay_pipe[4];
        int_delay_pipe[6]   <= int_delay_pipe[5];
        int_delay_pipe[7]   <= int_delay_pipe[6];
        int_delay_pipe[8]   <= int_delay_pipe[7];
        int_delay_pipe[9]   <= int_delay_pipe[8];
        int_delay_pipe[10]  <= int_delay_pipe[9];
        int_delay_pipe[11]  <= int_delay_pipe[10];
        int_delay_pipe[12]  <= int_delay_pipe[11];
        int_delay_pipe[13]  <= int_delay_pipe[12];
        int_delay_pipe[14]  <= int_delay_pipe[13];
        int_delay_pipe[15]  <= int_delay_pipe[14];
        int_delay_pipe[16]  <= int_delay_pipe[15];
        int_delay_pipe[17]  <= int_delay_pipe[16];
        int_delay_pipe[18]  <= int_delay_pipe[17];
        int_delay_pipe[19]  <= int_delay_pipe[18];
        int_delay_pipe[20]  <= int_delay_pipe[19];
        int_delay_pipe[21]  <= int_delay_pipe[20];
        int_delay_pipe[22]  <= int_delay_pipe[21];
        int_delay_pipe[23]  <= int_delay_pipe[22];
        int_delay_pipe[24]  <= int_delay_pipe[23];
        int_delay_pipe[25]  <= int_delay_pipe[24];
        int_delay_pipe[26]  <= int_delay_pipe[25];
        int_delay_pipe[27]  <= int_delay_pipe[26];
        int_delay_pipe[28]  <= int_delay_pipe[27];
        int_delay_pipe[29]  <= int_delay_pipe[28];
        int_delay_pipe[30]  <= int_delay_pipe[29];
        int_delay_pipe[31]  <= int_delay_pipe[30];
        int_delay_pipe[32]  <= int_delay_pipe[31];
        int_delay_pipe[33]  <= int_delay_pipe[32];
        int_delay_pipe[34]  <= int_delay_pipe[33];
        int_delay_pipe[35]  <= int_delay_pipe[34];
        int_delay_pipe[36]  <= int_delay_pipe[35];
        int_delay_pipe[37]  <= int_delay_pipe[36];
        int_delay_pipe[38]  <= int_delay_pipe[37];
        int_delay_pipe[39]  <= int_delay_pipe[38];
        int_delay_pipe[40]  <= int_delay_pipe[39];
        int_delay_pipe[41]  <= int_delay_pipe[40];
        int_delay_pipe[42]  <= int_delay_pipe[41];
        int_delay_pipe[43]  <= int_delay_pipe[42];
        int_delay_pipe[44]  <= int_delay_pipe[43];
        int_delay_pipe[45]  <= int_delay_pipe[44];
        int_delay_pipe[46]  <= int_delay_pipe[45];
        int_delay_pipe[47]  <= int_delay_pipe[46];
        int_delay_pipe[48]  <= int_delay_pipe[47];
        int_delay_pipe[49]  <= int_delay_pipe[48];
        int_delay_pipe[50]  <= int_delay_pipe[49];
        int_delay_pipe[51]  <= int_delay_pipe[50];
        int_delay_pipe[52]  <= int_delay_pipe[51];
        int_delay_pipe[53]  <= int_delay_pipe[52];
        int_delay_pipe[54]  <= int_delay_pipe[53];
        int_delay_pipe[55]  <= int_delay_pipe[54];
        int_delay_pipe[56]  <= int_delay_pipe[55];
        int_delay_pipe[57]  <= int_delay_pipe[56];
        int_delay_pipe[58]  <= int_delay_pipe[57];
        int_delay_pipe[59]  <= int_delay_pipe[58];
        int_delay_pipe[60]  <= int_delay_pipe[59];
        int_delay_pipe[61]  <= int_delay_pipe[60];
        int_delay_pipe[62]  <= int_delay_pipe[61];
        int_delay_pipe[63]  <= int_delay_pipe[62];
        int_delay_pipe[64]  <= int_delay_pipe[63];
        int_delay_pipe[65]  <= int_delay_pipe[64];
        int_delay_pipe[66]  <= int_delay_pipe[65];
        int_delay_pipe[67]  <= int_delay_pipe[66];
        int_delay_pipe[68]  <= int_delay_pipe[67];
        int_delay_pipe[69]  <= int_delay_pipe[68];
        int_delay_pipe[70]  <= int_delay_pipe[69];
        int_delay_pipe[71]  <= int_delay_pipe[70];
        int_delay_pipe[72]  <= int_delay_pipe[71];
        int_delay_pipe[73]  <= int_delay_pipe[72];
        int_delay_pipe[74]  <= int_delay_pipe[73];
        int_delay_pipe[75]  <= int_delay_pipe[74];
        int_delay_pipe[76]  <= int_delay_pipe[75];
        int_delay_pipe[77]  <= int_delay_pipe[76];
        int_delay_pipe[78]  <= int_delay_pipe[77];
        int_delay_pipe[79]  <= int_delay_pipe[78];
        int_delay_pipe[80]  <= int_delay_pipe[79];
        int_delay_pipe[81]  <= int_delay_pipe[80];
        int_delay_pipe[82]  <= int_delay_pipe[81];
        int_delay_pipe[83]  <= int_delay_pipe[82];
        int_delay_pipe[84]  <= int_delay_pipe[83];
        int_delay_pipe[85]  <= int_delay_pipe[84];
        int_delay_pipe[86]  <= int_delay_pipe[85];
        int_delay_pipe[87]  <= int_delay_pipe[86];
        int_delay_pipe[88]  <= int_delay_pipe[87];
        int_delay_pipe[89]  <= int_delay_pipe[88];
        int_delay_pipe[90]  <= int_delay_pipe[89];
        int_delay_pipe[91]  <= int_delay_pipe[90];
        int_delay_pipe[92]  <= int_delay_pipe[91];
        int_delay_pipe[93]  <= int_delay_pipe[92];
        int_delay_pipe[94]  <= int_delay_pipe[93];
        int_delay_pipe[95]  <= int_delay_pipe[94];
        int_delay_pipe[96]  <= int_delay_pipe[95];
        int_delay_pipe[97]  <= int_delay_pipe[96];
        int_delay_pipe[98]  <= int_delay_pipe[97];
        int_delay_pipe[99]  <= int_delay_pipe[98];
        int_delay_pipe[100] <= int_delay_pipe[99];
        int_delay_pipe[101] <= int_delay_pipe[100];
        int_delay_pipe[102] <= int_delay_pipe[101];
        int_delay_pipe[103] <= int_delay_pipe[102];
        int_delay_pipe[104] <= int_delay_pipe[103];
        int_delay_pipe[105] <= int_delay_pipe[104];
        int_delay_pipe[106] <= int_delay_pipe[105];
        int_delay_pipe[107] <= int_delay_pipe[106];
        int_delay_pipe[108] <= int_delay_pipe[107];
        int_delay_pipe[109] <= int_delay_pipe[108];
        int_delay_pipe[110] <= int_delay_pipe[109];
        int_delay_pipe[111] <= int_delay_pipe[110];
        int_delay_pipe[112] <= int_delay_pipe[111];
        int_delay_pipe[113] <= int_delay_pipe[112];
        int_delay_pipe[114] <= int_delay_pipe[113];
        int_delay_pipe[115] <= int_delay_pipe[114];
        int_delay_pipe[116] <= int_delay_pipe[115];
        int_delay_pipe[117] <= int_delay_pipe[116];
        int_delay_pipe[118] <= int_delay_pipe[117];
        int_delay_pipe[119] <= int_delay_pipe[118];
        int_delay_pipe[120] <= int_delay_pipe[119];
        int_delay_pipe[121] <= int_delay_pipe[120];
        int_delay_pipe[122] <= int_delay_pipe[121];
        int_delay_pipe[123] <= int_delay_pipe[122];
        int_delay_pipe[124] <= int_delay_pipe[123];
        int_delay_pipe[125] <= int_delay_pipe[124];
        int_delay_pipe[126] <= int_delay_pipe[125];
        int_delay_pipe[127] <= int_delay_pipe[126];
        int_delay_pipe[128] <= int_delay_pipe[127];
      end
    end
  end  // ceout_delayLine

  assign delayLine_out   = int_delay_pipe[128];

  assign expected_ce_out = delayLine_out & clk_enable;

  // -------------------------------------------------------------
  //  Checker: Checking the data received from the DUT.
  // -------------------------------------------------------------

  always @(posedge clk or posedge rst) begin
    filter_out_task(clk, rst, filter_out_rdenb, filter_out_addr, filter_out_done);
  end

  assign filter_out_rdenb = expected_ce_out;

  assign #clk_hold filter_out_dataTable = filter_out_expected[filter_out_addr];

  // ---- Bypass Register ----
  always @(posedge clk or posedge rst) begin : DataHoldRegister_temp_process2
    if (rst == 1'b1) begin
      regout <= 0;
    end else begin
      if (expected_ce_out == 1'b1) begin
        regout <= filter_out_dataTable;
      end
    end
  end  // DataHoldRegister_temp_process2

  assign filter_out_refTmp = (expected_ce_out == 1'b1) ? filter_out_dataTable : regout;


  assign filter_out_ref = filter_out_refTmp;



  always @ (posedge clk or posedge rst) // checker_filter_out
  begin
    if (rst == 1) begin
      filter_out_testFailure <= 0;
      filter_out_errCnt <= 0;
    end else begin
      if (filter_out_rdenb == 1) begin
        if (((abs(filter_out - filter_out_expected[filter_out_addr]) > 15) !== 0)) begin
          filter_out_errCnt <= filter_out_errCnt + 1;
          filter_out_testFailure <= 1;
          $display("ERROR  in filter_out at time %t : Expected '%h' Actual '%h'", $time,
                   filter_out_expected[filter_out_addr], filter_out);
          if (filter_out_errCnt >= MAX_ERROR_COUNT)
            $display(
                "Warning: Number of errors for filter_out have exceeded the maximum error limit"
            );
        end

      end
    end
  end  // checker_filter_out

  always @ (posedge clk or posedge rst) // checkDone_1
  begin
    if (rst == 1) check1_Done <= 0;
    else if ((check1_Done == 0) && (filter_out_done == 1) && (filter_out_rdenb == 1))
      check1_Done <= 1;
  end

  // -------------------------------------------------------------
  // Create done and test failure signal for output data
  // -------------------------------------------------------------

  assign snkDone = check1_Done;

  assign testFailure = filter_out_testFailure;

  // -------------------------------------------------------------
  // Global clock enable
  // -------------------------------------------------------------
  always @(snkDone, tbenb_dly) begin
    if (snkDone == 0) #clk_hold clk_enable <= tbenb_dly;
    else #clk_hold clk_enable <= 0;
  end

  // Assignment Statements



endmodule  // filter_impluse_tb
